// IMPORTANT NOTE: if using VPR, any instantiated BELs with no outputs MUST be instantiated after IO
// This is because VPR auto-generates names for primitives with no outputs, and we assume OutPass BELs
// are the first BELs to be auto-named in our constraints file.

module template ();
wire Tile_X0Y1_A_I, Tile_X0Y1_A_T, Tile_X0Y1_A_O, Tile_X0Y1_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y1_A (.O(Tile_X0Y1_A_O), .Q(Tile_X0Y1_A_Q), .I(Tile_X0Y1_A_I));

wire Tile_X0Y1_B_I, Tile_X0Y1_B_T, Tile_X0Y1_B_O, Tile_X0Y1_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y1_B (.O(Tile_X0Y1_B_O), .Q(Tile_X0Y1_B_Q), .I(Tile_X0Y1_B_I));

wire Tile_X10Y1_RAM2FAB_D0_O0, Tile_X10Y1_RAM2FAB_D0_O1, Tile_X10Y1_RAM2FAB_D0_O2, Tile_X10Y1_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X10Y1_A (.O0(Tile_X10Y1_RAM2FAB_D0_O0), .O1(Tile_X10Y1_RAM2FAB_D0_O1), .O2(Tile_X10Y1_RAM2FAB_D0_O2), .O3(Tile_X10Y1_RAM2FAB_D0_O3));

wire Tile_X10Y1_RAM2FAB_D1_O0, Tile_X10Y1_RAM2FAB_D1_O1, Tile_X10Y1_RAM2FAB_D1_O2, Tile_X10Y1_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X10Y1_B (.O0(Tile_X10Y1_RAM2FAB_D1_O0), .O1(Tile_X10Y1_RAM2FAB_D1_O1), .O2(Tile_X10Y1_RAM2FAB_D1_O2), .O3(Tile_X10Y1_RAM2FAB_D1_O3));

wire Tile_X10Y1_RAM2FAB_D2_O0, Tile_X10Y1_RAM2FAB_D2_O1, Tile_X10Y1_RAM2FAB_D2_O2, Tile_X10Y1_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X10Y1_C (.O0(Tile_X10Y1_RAM2FAB_D2_O0), .O1(Tile_X10Y1_RAM2FAB_D2_O1), .O2(Tile_X10Y1_RAM2FAB_D2_O2), .O3(Tile_X10Y1_RAM2FAB_D2_O3));

wire Tile_X10Y1_RAM2FAB_D3_O0, Tile_X10Y1_RAM2FAB_D3_O1, Tile_X10Y1_RAM2FAB_D3_O2, Tile_X10Y1_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X10Y1_D (.O0(Tile_X10Y1_RAM2FAB_D3_O0), .O1(Tile_X10Y1_RAM2FAB_D3_O1), .O2(Tile_X10Y1_RAM2FAB_D3_O2), .O3(Tile_X10Y1_RAM2FAB_D3_O3));

wire Tile_X10Y1_FAB2RAM_D0_I0, Tile_X10Y1_FAB2RAM_D0_I1, Tile_X10Y1_FAB2RAM_D0_I2, Tile_X10Y1_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y1_E (.I0(Tile_X10Y1_FAB2RAM_D0_I0), .I1(Tile_X10Y1_FAB2RAM_D0_I1), .I2(Tile_X10Y1_FAB2RAM_D0_I2), .I3(Tile_X10Y1_FAB2RAM_D0_I3));

wire Tile_X10Y1_FAB2RAM_D1_I0, Tile_X10Y1_FAB2RAM_D1_I1, Tile_X10Y1_FAB2RAM_D1_I2, Tile_X10Y1_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y1_F (.I0(Tile_X10Y1_FAB2RAM_D1_I0), .I1(Tile_X10Y1_FAB2RAM_D1_I1), .I2(Tile_X10Y1_FAB2RAM_D1_I2), .I3(Tile_X10Y1_FAB2RAM_D1_I3));

wire Tile_X10Y1_FAB2RAM_D2_I0, Tile_X10Y1_FAB2RAM_D2_I1, Tile_X10Y1_FAB2RAM_D2_I2, Tile_X10Y1_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X10Y1_G (.I0(Tile_X10Y1_FAB2RAM_D2_I0), .I1(Tile_X10Y1_FAB2RAM_D2_I1), .I2(Tile_X10Y1_FAB2RAM_D2_I2), .I3(Tile_X10Y1_FAB2RAM_D2_I3));

wire Tile_X10Y1_FAB2RAM_D3_I0, Tile_X10Y1_FAB2RAM_D3_I1, Tile_X10Y1_FAB2RAM_D3_I2, Tile_X10Y1_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X10Y1_H (.I0(Tile_X10Y1_FAB2RAM_D3_I0), .I1(Tile_X10Y1_FAB2RAM_D3_I1), .I2(Tile_X10Y1_FAB2RAM_D3_I2), .I3(Tile_X10Y1_FAB2RAM_D3_I3));

wire Tile_X10Y1_FAB2RAM_A0_I0, Tile_X10Y1_FAB2RAM_A0_I1, Tile_X10Y1_FAB2RAM_A0_I2, Tile_X10Y1_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y1_I (.I0(Tile_X10Y1_FAB2RAM_A0_I0), .I1(Tile_X10Y1_FAB2RAM_A0_I1), .I2(Tile_X10Y1_FAB2RAM_A0_I2), .I3(Tile_X10Y1_FAB2RAM_A0_I3));

wire Tile_X10Y1_FAB2RAM_A1_I0, Tile_X10Y1_FAB2RAM_A1_I1, Tile_X10Y1_FAB2RAM_A1_I2, Tile_X10Y1_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y1_J (.I0(Tile_X10Y1_FAB2RAM_A1_I0), .I1(Tile_X10Y1_FAB2RAM_A1_I1), .I2(Tile_X10Y1_FAB2RAM_A1_I2), .I3(Tile_X10Y1_FAB2RAM_A1_I3));

wire Tile_X10Y1_FAB2RAM_C_I0, Tile_X10Y1_FAB2RAM_C_I1, Tile_X10Y1_FAB2RAM_C_I2, Tile_X10Y1_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X10Y1_K (.I0(Tile_X10Y1_FAB2RAM_C_I0), .I1(Tile_X10Y1_FAB2RAM_C_I1), .I2(Tile_X10Y1_FAB2RAM_C_I2), .I3(Tile_X10Y1_FAB2RAM_C_I3));

wire Tile_X0Y2_A_I, Tile_X0Y2_A_T, Tile_X0Y2_A_O, Tile_X0Y2_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y2_A (.O(Tile_X0Y2_A_O), .Q(Tile_X0Y2_A_Q), .I(Tile_X0Y2_A_I));

wire Tile_X0Y2_B_I, Tile_X0Y2_B_T, Tile_X0Y2_B_O, Tile_X0Y2_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y2_B (.O(Tile_X0Y2_B_O), .Q(Tile_X0Y2_B_Q), .I(Tile_X0Y2_B_I));

wire Tile_X10Y2_RAM2FAB_D0_O0, Tile_X10Y2_RAM2FAB_D0_O1, Tile_X10Y2_RAM2FAB_D0_O2, Tile_X10Y2_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X10Y2_A (.O0(Tile_X10Y2_RAM2FAB_D0_O0), .O1(Tile_X10Y2_RAM2FAB_D0_O1), .O2(Tile_X10Y2_RAM2FAB_D0_O2), .O3(Tile_X10Y2_RAM2FAB_D0_O3));

wire Tile_X10Y2_RAM2FAB_D1_O0, Tile_X10Y2_RAM2FAB_D1_O1, Tile_X10Y2_RAM2FAB_D1_O2, Tile_X10Y2_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X10Y2_B (.O0(Tile_X10Y2_RAM2FAB_D1_O0), .O1(Tile_X10Y2_RAM2FAB_D1_O1), .O2(Tile_X10Y2_RAM2FAB_D1_O2), .O3(Tile_X10Y2_RAM2FAB_D1_O3));

wire Tile_X10Y2_RAM2FAB_D2_O0, Tile_X10Y2_RAM2FAB_D2_O1, Tile_X10Y2_RAM2FAB_D2_O2, Tile_X10Y2_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X10Y2_C (.O0(Tile_X10Y2_RAM2FAB_D2_O0), .O1(Tile_X10Y2_RAM2FAB_D2_O1), .O2(Tile_X10Y2_RAM2FAB_D2_O2), .O3(Tile_X10Y2_RAM2FAB_D2_O3));

wire Tile_X10Y2_RAM2FAB_D3_O0, Tile_X10Y2_RAM2FAB_D3_O1, Tile_X10Y2_RAM2FAB_D3_O2, Tile_X10Y2_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X10Y2_D (.O0(Tile_X10Y2_RAM2FAB_D3_O0), .O1(Tile_X10Y2_RAM2FAB_D3_O1), .O2(Tile_X10Y2_RAM2FAB_D3_O2), .O3(Tile_X10Y2_RAM2FAB_D3_O3));

wire Tile_X10Y2_FAB2RAM_D0_I0, Tile_X10Y2_FAB2RAM_D0_I1, Tile_X10Y2_FAB2RAM_D0_I2, Tile_X10Y2_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y2_E (.I0(Tile_X10Y2_FAB2RAM_D0_I0), .I1(Tile_X10Y2_FAB2RAM_D0_I1), .I2(Tile_X10Y2_FAB2RAM_D0_I2), .I3(Tile_X10Y2_FAB2RAM_D0_I3));

wire Tile_X10Y2_FAB2RAM_D1_I0, Tile_X10Y2_FAB2RAM_D1_I1, Tile_X10Y2_FAB2RAM_D1_I2, Tile_X10Y2_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y2_F (.I0(Tile_X10Y2_FAB2RAM_D1_I0), .I1(Tile_X10Y2_FAB2RAM_D1_I1), .I2(Tile_X10Y2_FAB2RAM_D1_I2), .I3(Tile_X10Y2_FAB2RAM_D1_I3));

wire Tile_X10Y2_FAB2RAM_D2_I0, Tile_X10Y2_FAB2RAM_D2_I1, Tile_X10Y2_FAB2RAM_D2_I2, Tile_X10Y2_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X10Y2_G (.I0(Tile_X10Y2_FAB2RAM_D2_I0), .I1(Tile_X10Y2_FAB2RAM_D2_I1), .I2(Tile_X10Y2_FAB2RAM_D2_I2), .I3(Tile_X10Y2_FAB2RAM_D2_I3));

wire Tile_X10Y2_FAB2RAM_D3_I0, Tile_X10Y2_FAB2RAM_D3_I1, Tile_X10Y2_FAB2RAM_D3_I2, Tile_X10Y2_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X10Y2_H (.I0(Tile_X10Y2_FAB2RAM_D3_I0), .I1(Tile_X10Y2_FAB2RAM_D3_I1), .I2(Tile_X10Y2_FAB2RAM_D3_I2), .I3(Tile_X10Y2_FAB2RAM_D3_I3));

wire Tile_X10Y2_FAB2RAM_A0_I0, Tile_X10Y2_FAB2RAM_A0_I1, Tile_X10Y2_FAB2RAM_A0_I2, Tile_X10Y2_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y2_I (.I0(Tile_X10Y2_FAB2RAM_A0_I0), .I1(Tile_X10Y2_FAB2RAM_A0_I1), .I2(Tile_X10Y2_FAB2RAM_A0_I2), .I3(Tile_X10Y2_FAB2RAM_A0_I3));

wire Tile_X10Y2_FAB2RAM_A1_I0, Tile_X10Y2_FAB2RAM_A1_I1, Tile_X10Y2_FAB2RAM_A1_I2, Tile_X10Y2_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y2_J (.I0(Tile_X10Y2_FAB2RAM_A1_I0), .I1(Tile_X10Y2_FAB2RAM_A1_I1), .I2(Tile_X10Y2_FAB2RAM_A1_I2), .I3(Tile_X10Y2_FAB2RAM_A1_I3));

wire Tile_X10Y2_FAB2RAM_C_I0, Tile_X10Y2_FAB2RAM_C_I1, Tile_X10Y2_FAB2RAM_C_I2, Tile_X10Y2_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X10Y2_K (.I0(Tile_X10Y2_FAB2RAM_C_I0), .I1(Tile_X10Y2_FAB2RAM_C_I1), .I2(Tile_X10Y2_FAB2RAM_C_I2), .I3(Tile_X10Y2_FAB2RAM_C_I3));

wire Tile_X0Y3_A_I, Tile_X0Y3_A_T, Tile_X0Y3_A_O, Tile_X0Y3_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y3_A (.O(Tile_X0Y3_A_O), .Q(Tile_X0Y3_A_Q), .I(Tile_X0Y3_A_I));

wire Tile_X0Y3_B_I, Tile_X0Y3_B_T, Tile_X0Y3_B_O, Tile_X0Y3_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y3_B (.O(Tile_X0Y3_B_O), .Q(Tile_X0Y3_B_Q), .I(Tile_X0Y3_B_I));

wire Tile_X10Y3_RAM2FAB_D0_O0, Tile_X10Y3_RAM2FAB_D0_O1, Tile_X10Y3_RAM2FAB_D0_O2, Tile_X10Y3_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X10Y3_A (.O0(Tile_X10Y3_RAM2FAB_D0_O0), .O1(Tile_X10Y3_RAM2FAB_D0_O1), .O2(Tile_X10Y3_RAM2FAB_D0_O2), .O3(Tile_X10Y3_RAM2FAB_D0_O3));

wire Tile_X10Y3_RAM2FAB_D1_O0, Tile_X10Y3_RAM2FAB_D1_O1, Tile_X10Y3_RAM2FAB_D1_O2, Tile_X10Y3_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X10Y3_B (.O0(Tile_X10Y3_RAM2FAB_D1_O0), .O1(Tile_X10Y3_RAM2FAB_D1_O1), .O2(Tile_X10Y3_RAM2FAB_D1_O2), .O3(Tile_X10Y3_RAM2FAB_D1_O3));

wire Tile_X10Y3_RAM2FAB_D2_O0, Tile_X10Y3_RAM2FAB_D2_O1, Tile_X10Y3_RAM2FAB_D2_O2, Tile_X10Y3_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X10Y3_C (.O0(Tile_X10Y3_RAM2FAB_D2_O0), .O1(Tile_X10Y3_RAM2FAB_D2_O1), .O2(Tile_X10Y3_RAM2FAB_D2_O2), .O3(Tile_X10Y3_RAM2FAB_D2_O3));

wire Tile_X10Y3_RAM2FAB_D3_O0, Tile_X10Y3_RAM2FAB_D3_O1, Tile_X10Y3_RAM2FAB_D3_O2, Tile_X10Y3_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X10Y3_D (.O0(Tile_X10Y3_RAM2FAB_D3_O0), .O1(Tile_X10Y3_RAM2FAB_D3_O1), .O2(Tile_X10Y3_RAM2FAB_D3_O2), .O3(Tile_X10Y3_RAM2FAB_D3_O3));

wire Tile_X10Y3_FAB2RAM_D0_I0, Tile_X10Y3_FAB2RAM_D0_I1, Tile_X10Y3_FAB2RAM_D0_I2, Tile_X10Y3_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y3_E (.I0(Tile_X10Y3_FAB2RAM_D0_I0), .I1(Tile_X10Y3_FAB2RAM_D0_I1), .I2(Tile_X10Y3_FAB2RAM_D0_I2), .I3(Tile_X10Y3_FAB2RAM_D0_I3));

wire Tile_X10Y3_FAB2RAM_D1_I0, Tile_X10Y3_FAB2RAM_D1_I1, Tile_X10Y3_FAB2RAM_D1_I2, Tile_X10Y3_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y3_F (.I0(Tile_X10Y3_FAB2RAM_D1_I0), .I1(Tile_X10Y3_FAB2RAM_D1_I1), .I2(Tile_X10Y3_FAB2RAM_D1_I2), .I3(Tile_X10Y3_FAB2RAM_D1_I3));

wire Tile_X10Y3_FAB2RAM_D2_I0, Tile_X10Y3_FAB2RAM_D2_I1, Tile_X10Y3_FAB2RAM_D2_I2, Tile_X10Y3_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X10Y3_G (.I0(Tile_X10Y3_FAB2RAM_D2_I0), .I1(Tile_X10Y3_FAB2RAM_D2_I1), .I2(Tile_X10Y3_FAB2RAM_D2_I2), .I3(Tile_X10Y3_FAB2RAM_D2_I3));

wire Tile_X10Y3_FAB2RAM_D3_I0, Tile_X10Y3_FAB2RAM_D3_I1, Tile_X10Y3_FAB2RAM_D3_I2, Tile_X10Y3_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X10Y3_H (.I0(Tile_X10Y3_FAB2RAM_D3_I0), .I1(Tile_X10Y3_FAB2RAM_D3_I1), .I2(Tile_X10Y3_FAB2RAM_D3_I2), .I3(Tile_X10Y3_FAB2RAM_D3_I3));

wire Tile_X10Y3_FAB2RAM_A0_I0, Tile_X10Y3_FAB2RAM_A0_I1, Tile_X10Y3_FAB2RAM_A0_I2, Tile_X10Y3_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y3_I (.I0(Tile_X10Y3_FAB2RAM_A0_I0), .I1(Tile_X10Y3_FAB2RAM_A0_I1), .I2(Tile_X10Y3_FAB2RAM_A0_I2), .I3(Tile_X10Y3_FAB2RAM_A0_I3));

wire Tile_X10Y3_FAB2RAM_A1_I0, Tile_X10Y3_FAB2RAM_A1_I1, Tile_X10Y3_FAB2RAM_A1_I2, Tile_X10Y3_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y3_J (.I0(Tile_X10Y3_FAB2RAM_A1_I0), .I1(Tile_X10Y3_FAB2RAM_A1_I1), .I2(Tile_X10Y3_FAB2RAM_A1_I2), .I3(Tile_X10Y3_FAB2RAM_A1_I3));

wire Tile_X10Y3_FAB2RAM_C_I0, Tile_X10Y3_FAB2RAM_C_I1, Tile_X10Y3_FAB2RAM_C_I2, Tile_X10Y3_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X10Y3_K (.I0(Tile_X10Y3_FAB2RAM_C_I0), .I1(Tile_X10Y3_FAB2RAM_C_I1), .I2(Tile_X10Y3_FAB2RAM_C_I2), .I3(Tile_X10Y3_FAB2RAM_C_I3));

wire Tile_X0Y4_A_I, Tile_X0Y4_A_T, Tile_X0Y4_A_O, Tile_X0Y4_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y4_A (.O(Tile_X0Y4_A_O), .Q(Tile_X0Y4_A_Q), .I(Tile_X0Y4_A_I));

wire Tile_X0Y4_B_I, Tile_X0Y4_B_T, Tile_X0Y4_B_O, Tile_X0Y4_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y4_B (.O(Tile_X0Y4_B_O), .Q(Tile_X0Y4_B_Q), .I(Tile_X0Y4_B_I));

wire Tile_X10Y4_RAM2FAB_D0_O0, Tile_X10Y4_RAM2FAB_D0_O1, Tile_X10Y4_RAM2FAB_D0_O2, Tile_X10Y4_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X10Y4_A (.O0(Tile_X10Y4_RAM2FAB_D0_O0), .O1(Tile_X10Y4_RAM2FAB_D0_O1), .O2(Tile_X10Y4_RAM2FAB_D0_O2), .O3(Tile_X10Y4_RAM2FAB_D0_O3));

wire Tile_X10Y4_RAM2FAB_D1_O0, Tile_X10Y4_RAM2FAB_D1_O1, Tile_X10Y4_RAM2FAB_D1_O2, Tile_X10Y4_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X10Y4_B (.O0(Tile_X10Y4_RAM2FAB_D1_O0), .O1(Tile_X10Y4_RAM2FAB_D1_O1), .O2(Tile_X10Y4_RAM2FAB_D1_O2), .O3(Tile_X10Y4_RAM2FAB_D1_O3));

wire Tile_X10Y4_RAM2FAB_D2_O0, Tile_X10Y4_RAM2FAB_D2_O1, Tile_X10Y4_RAM2FAB_D2_O2, Tile_X10Y4_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X10Y4_C (.O0(Tile_X10Y4_RAM2FAB_D2_O0), .O1(Tile_X10Y4_RAM2FAB_D2_O1), .O2(Tile_X10Y4_RAM2FAB_D2_O2), .O3(Tile_X10Y4_RAM2FAB_D2_O3));

wire Tile_X10Y4_RAM2FAB_D3_O0, Tile_X10Y4_RAM2FAB_D3_O1, Tile_X10Y4_RAM2FAB_D3_O2, Tile_X10Y4_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X10Y4_D (.O0(Tile_X10Y4_RAM2FAB_D3_O0), .O1(Tile_X10Y4_RAM2FAB_D3_O1), .O2(Tile_X10Y4_RAM2FAB_D3_O2), .O3(Tile_X10Y4_RAM2FAB_D3_O3));

wire Tile_X10Y4_FAB2RAM_D0_I0, Tile_X10Y4_FAB2RAM_D0_I1, Tile_X10Y4_FAB2RAM_D0_I2, Tile_X10Y4_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y4_E (.I0(Tile_X10Y4_FAB2RAM_D0_I0), .I1(Tile_X10Y4_FAB2RAM_D0_I1), .I2(Tile_X10Y4_FAB2RAM_D0_I2), .I3(Tile_X10Y4_FAB2RAM_D0_I3));

wire Tile_X10Y4_FAB2RAM_D1_I0, Tile_X10Y4_FAB2RAM_D1_I1, Tile_X10Y4_FAB2RAM_D1_I2, Tile_X10Y4_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y4_F (.I0(Tile_X10Y4_FAB2RAM_D1_I0), .I1(Tile_X10Y4_FAB2RAM_D1_I1), .I2(Tile_X10Y4_FAB2RAM_D1_I2), .I3(Tile_X10Y4_FAB2RAM_D1_I3));

wire Tile_X10Y4_FAB2RAM_D2_I0, Tile_X10Y4_FAB2RAM_D2_I1, Tile_X10Y4_FAB2RAM_D2_I2, Tile_X10Y4_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X10Y4_G (.I0(Tile_X10Y4_FAB2RAM_D2_I0), .I1(Tile_X10Y4_FAB2RAM_D2_I1), .I2(Tile_X10Y4_FAB2RAM_D2_I2), .I3(Tile_X10Y4_FAB2RAM_D2_I3));

wire Tile_X10Y4_FAB2RAM_D3_I0, Tile_X10Y4_FAB2RAM_D3_I1, Tile_X10Y4_FAB2RAM_D3_I2, Tile_X10Y4_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X10Y4_H (.I0(Tile_X10Y4_FAB2RAM_D3_I0), .I1(Tile_X10Y4_FAB2RAM_D3_I1), .I2(Tile_X10Y4_FAB2RAM_D3_I2), .I3(Tile_X10Y4_FAB2RAM_D3_I3));

wire Tile_X10Y4_FAB2RAM_A0_I0, Tile_X10Y4_FAB2RAM_A0_I1, Tile_X10Y4_FAB2RAM_A0_I2, Tile_X10Y4_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y4_I (.I0(Tile_X10Y4_FAB2RAM_A0_I0), .I1(Tile_X10Y4_FAB2RAM_A0_I1), .I2(Tile_X10Y4_FAB2RAM_A0_I2), .I3(Tile_X10Y4_FAB2RAM_A0_I3));

wire Tile_X10Y4_FAB2RAM_A1_I0, Tile_X10Y4_FAB2RAM_A1_I1, Tile_X10Y4_FAB2RAM_A1_I2, Tile_X10Y4_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y4_J (.I0(Tile_X10Y4_FAB2RAM_A1_I0), .I1(Tile_X10Y4_FAB2RAM_A1_I1), .I2(Tile_X10Y4_FAB2RAM_A1_I2), .I3(Tile_X10Y4_FAB2RAM_A1_I3));

wire Tile_X10Y4_FAB2RAM_C_I0, Tile_X10Y4_FAB2RAM_C_I1, Tile_X10Y4_FAB2RAM_C_I2, Tile_X10Y4_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X10Y4_K (.I0(Tile_X10Y4_FAB2RAM_C_I0), .I1(Tile_X10Y4_FAB2RAM_C_I1), .I2(Tile_X10Y4_FAB2RAM_C_I2), .I3(Tile_X10Y4_FAB2RAM_C_I3));

wire Tile_X0Y5_A_I, Tile_X0Y5_A_T, Tile_X0Y5_A_O, Tile_X0Y5_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y5_A (.O(Tile_X0Y5_A_O), .Q(Tile_X0Y5_A_Q), .I(Tile_X0Y5_A_I));

wire Tile_X0Y5_B_I, Tile_X0Y5_B_T, Tile_X0Y5_B_O, Tile_X0Y5_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y5_B (.O(Tile_X0Y5_B_O), .Q(Tile_X0Y5_B_Q), .I(Tile_X0Y5_B_I));

wire Tile_X10Y5_RAM2FAB_D0_O0, Tile_X10Y5_RAM2FAB_D0_O1, Tile_X10Y5_RAM2FAB_D0_O2, Tile_X10Y5_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X10Y5_A (.O0(Tile_X10Y5_RAM2FAB_D0_O0), .O1(Tile_X10Y5_RAM2FAB_D0_O1), .O2(Tile_X10Y5_RAM2FAB_D0_O2), .O3(Tile_X10Y5_RAM2FAB_D0_O3));

wire Tile_X10Y5_RAM2FAB_D1_O0, Tile_X10Y5_RAM2FAB_D1_O1, Tile_X10Y5_RAM2FAB_D1_O2, Tile_X10Y5_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X10Y5_B (.O0(Tile_X10Y5_RAM2FAB_D1_O0), .O1(Tile_X10Y5_RAM2FAB_D1_O1), .O2(Tile_X10Y5_RAM2FAB_D1_O2), .O3(Tile_X10Y5_RAM2FAB_D1_O3));

wire Tile_X10Y5_RAM2FAB_D2_O0, Tile_X10Y5_RAM2FAB_D2_O1, Tile_X10Y5_RAM2FAB_D2_O2, Tile_X10Y5_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X10Y5_C (.O0(Tile_X10Y5_RAM2FAB_D2_O0), .O1(Tile_X10Y5_RAM2FAB_D2_O1), .O2(Tile_X10Y5_RAM2FAB_D2_O2), .O3(Tile_X10Y5_RAM2FAB_D2_O3));

wire Tile_X10Y5_RAM2FAB_D3_O0, Tile_X10Y5_RAM2FAB_D3_O1, Tile_X10Y5_RAM2FAB_D3_O2, Tile_X10Y5_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X10Y5_D (.O0(Tile_X10Y5_RAM2FAB_D3_O0), .O1(Tile_X10Y5_RAM2FAB_D3_O1), .O2(Tile_X10Y5_RAM2FAB_D3_O2), .O3(Tile_X10Y5_RAM2FAB_D3_O3));

wire Tile_X10Y5_FAB2RAM_D0_I0, Tile_X10Y5_FAB2RAM_D0_I1, Tile_X10Y5_FAB2RAM_D0_I2, Tile_X10Y5_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y5_E (.I0(Tile_X10Y5_FAB2RAM_D0_I0), .I1(Tile_X10Y5_FAB2RAM_D0_I1), .I2(Tile_X10Y5_FAB2RAM_D0_I2), .I3(Tile_X10Y5_FAB2RAM_D0_I3));

wire Tile_X10Y5_FAB2RAM_D1_I0, Tile_X10Y5_FAB2RAM_D1_I1, Tile_X10Y5_FAB2RAM_D1_I2, Tile_X10Y5_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y5_F (.I0(Tile_X10Y5_FAB2RAM_D1_I0), .I1(Tile_X10Y5_FAB2RAM_D1_I1), .I2(Tile_X10Y5_FAB2RAM_D1_I2), .I3(Tile_X10Y5_FAB2RAM_D1_I3));

wire Tile_X10Y5_FAB2RAM_D2_I0, Tile_X10Y5_FAB2RAM_D2_I1, Tile_X10Y5_FAB2RAM_D2_I2, Tile_X10Y5_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X10Y5_G (.I0(Tile_X10Y5_FAB2RAM_D2_I0), .I1(Tile_X10Y5_FAB2RAM_D2_I1), .I2(Tile_X10Y5_FAB2RAM_D2_I2), .I3(Tile_X10Y5_FAB2RAM_D2_I3));

wire Tile_X10Y5_FAB2RAM_D3_I0, Tile_X10Y5_FAB2RAM_D3_I1, Tile_X10Y5_FAB2RAM_D3_I2, Tile_X10Y5_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X10Y5_H (.I0(Tile_X10Y5_FAB2RAM_D3_I0), .I1(Tile_X10Y5_FAB2RAM_D3_I1), .I2(Tile_X10Y5_FAB2RAM_D3_I2), .I3(Tile_X10Y5_FAB2RAM_D3_I3));

wire Tile_X10Y5_FAB2RAM_A0_I0, Tile_X10Y5_FAB2RAM_A0_I1, Tile_X10Y5_FAB2RAM_A0_I2, Tile_X10Y5_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y5_I (.I0(Tile_X10Y5_FAB2RAM_A0_I0), .I1(Tile_X10Y5_FAB2RAM_A0_I1), .I2(Tile_X10Y5_FAB2RAM_A0_I2), .I3(Tile_X10Y5_FAB2RAM_A0_I3));

wire Tile_X10Y5_FAB2RAM_A1_I0, Tile_X10Y5_FAB2RAM_A1_I1, Tile_X10Y5_FAB2RAM_A1_I2, Tile_X10Y5_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y5_J (.I0(Tile_X10Y5_FAB2RAM_A1_I0), .I1(Tile_X10Y5_FAB2RAM_A1_I1), .I2(Tile_X10Y5_FAB2RAM_A1_I2), .I3(Tile_X10Y5_FAB2RAM_A1_I3));

wire Tile_X10Y5_FAB2RAM_C_I0, Tile_X10Y5_FAB2RAM_C_I1, Tile_X10Y5_FAB2RAM_C_I2, Tile_X10Y5_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X10Y5_K (.I0(Tile_X10Y5_FAB2RAM_C_I0), .I1(Tile_X10Y5_FAB2RAM_C_I1), .I2(Tile_X10Y5_FAB2RAM_C_I2), .I3(Tile_X10Y5_FAB2RAM_C_I3));

wire Tile_X0Y6_A_I, Tile_X0Y6_A_T, Tile_X0Y6_A_O, Tile_X0Y6_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y6_A (.O(Tile_X0Y6_A_O), .Q(Tile_X0Y6_A_Q), .I(Tile_X0Y6_A_I));

wire Tile_X0Y6_B_I, Tile_X0Y6_B_T, Tile_X0Y6_B_O, Tile_X0Y6_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y6_B (.O(Tile_X0Y6_B_O), .Q(Tile_X0Y6_B_Q), .I(Tile_X0Y6_B_I));

wire Tile_X10Y6_RAM2FAB_D0_O0, Tile_X10Y6_RAM2FAB_D0_O1, Tile_X10Y6_RAM2FAB_D0_O2, Tile_X10Y6_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X10Y6_A (.O0(Tile_X10Y6_RAM2FAB_D0_O0), .O1(Tile_X10Y6_RAM2FAB_D0_O1), .O2(Tile_X10Y6_RAM2FAB_D0_O2), .O3(Tile_X10Y6_RAM2FAB_D0_O3));

wire Tile_X10Y6_RAM2FAB_D1_O0, Tile_X10Y6_RAM2FAB_D1_O1, Tile_X10Y6_RAM2FAB_D1_O2, Tile_X10Y6_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X10Y6_B (.O0(Tile_X10Y6_RAM2FAB_D1_O0), .O1(Tile_X10Y6_RAM2FAB_D1_O1), .O2(Tile_X10Y6_RAM2FAB_D1_O2), .O3(Tile_X10Y6_RAM2FAB_D1_O3));

wire Tile_X10Y6_RAM2FAB_D2_O0, Tile_X10Y6_RAM2FAB_D2_O1, Tile_X10Y6_RAM2FAB_D2_O2, Tile_X10Y6_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X10Y6_C (.O0(Tile_X10Y6_RAM2FAB_D2_O0), .O1(Tile_X10Y6_RAM2FAB_D2_O1), .O2(Tile_X10Y6_RAM2FAB_D2_O2), .O3(Tile_X10Y6_RAM2FAB_D2_O3));

wire Tile_X10Y6_RAM2FAB_D3_O0, Tile_X10Y6_RAM2FAB_D3_O1, Tile_X10Y6_RAM2FAB_D3_O2, Tile_X10Y6_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X10Y6_D (.O0(Tile_X10Y6_RAM2FAB_D3_O0), .O1(Tile_X10Y6_RAM2FAB_D3_O1), .O2(Tile_X10Y6_RAM2FAB_D3_O2), .O3(Tile_X10Y6_RAM2FAB_D3_O3));

wire Tile_X10Y6_FAB2RAM_D0_I0, Tile_X10Y6_FAB2RAM_D0_I1, Tile_X10Y6_FAB2RAM_D0_I2, Tile_X10Y6_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y6_E (.I0(Tile_X10Y6_FAB2RAM_D0_I0), .I1(Tile_X10Y6_FAB2RAM_D0_I1), .I2(Tile_X10Y6_FAB2RAM_D0_I2), .I3(Tile_X10Y6_FAB2RAM_D0_I3));

wire Tile_X10Y6_FAB2RAM_D1_I0, Tile_X10Y6_FAB2RAM_D1_I1, Tile_X10Y6_FAB2RAM_D1_I2, Tile_X10Y6_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y6_F (.I0(Tile_X10Y6_FAB2RAM_D1_I0), .I1(Tile_X10Y6_FAB2RAM_D1_I1), .I2(Tile_X10Y6_FAB2RAM_D1_I2), .I3(Tile_X10Y6_FAB2RAM_D1_I3));

wire Tile_X10Y6_FAB2RAM_D2_I0, Tile_X10Y6_FAB2RAM_D2_I1, Tile_X10Y6_FAB2RAM_D2_I2, Tile_X10Y6_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X10Y6_G (.I0(Tile_X10Y6_FAB2RAM_D2_I0), .I1(Tile_X10Y6_FAB2RAM_D2_I1), .I2(Tile_X10Y6_FAB2RAM_D2_I2), .I3(Tile_X10Y6_FAB2RAM_D2_I3));

wire Tile_X10Y6_FAB2RAM_D3_I0, Tile_X10Y6_FAB2RAM_D3_I1, Tile_X10Y6_FAB2RAM_D3_I2, Tile_X10Y6_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X10Y6_H (.I0(Tile_X10Y6_FAB2RAM_D3_I0), .I1(Tile_X10Y6_FAB2RAM_D3_I1), .I2(Tile_X10Y6_FAB2RAM_D3_I2), .I3(Tile_X10Y6_FAB2RAM_D3_I3));

wire Tile_X10Y6_FAB2RAM_A0_I0, Tile_X10Y6_FAB2RAM_A0_I1, Tile_X10Y6_FAB2RAM_A0_I2, Tile_X10Y6_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y6_I (.I0(Tile_X10Y6_FAB2RAM_A0_I0), .I1(Tile_X10Y6_FAB2RAM_A0_I1), .I2(Tile_X10Y6_FAB2RAM_A0_I2), .I3(Tile_X10Y6_FAB2RAM_A0_I3));

wire Tile_X10Y6_FAB2RAM_A1_I0, Tile_X10Y6_FAB2RAM_A1_I1, Tile_X10Y6_FAB2RAM_A1_I2, Tile_X10Y6_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y6_J (.I0(Tile_X10Y6_FAB2RAM_A1_I0), .I1(Tile_X10Y6_FAB2RAM_A1_I1), .I2(Tile_X10Y6_FAB2RAM_A1_I2), .I3(Tile_X10Y6_FAB2RAM_A1_I3));

wire Tile_X10Y6_FAB2RAM_C_I0, Tile_X10Y6_FAB2RAM_C_I1, Tile_X10Y6_FAB2RAM_C_I2, Tile_X10Y6_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X10Y6_K (.I0(Tile_X10Y6_FAB2RAM_C_I0), .I1(Tile_X10Y6_FAB2RAM_C_I1), .I2(Tile_X10Y6_FAB2RAM_C_I2), .I3(Tile_X10Y6_FAB2RAM_C_I3));

wire Tile_X0Y7_A_I, Tile_X0Y7_A_T, Tile_X0Y7_A_O, Tile_X0Y7_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y7_A (.O(Tile_X0Y7_A_O), .Q(Tile_X0Y7_A_Q), .I(Tile_X0Y7_A_I));

wire Tile_X0Y7_B_I, Tile_X0Y7_B_T, Tile_X0Y7_B_O, Tile_X0Y7_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y7_B (.O(Tile_X0Y7_B_O), .Q(Tile_X0Y7_B_Q), .I(Tile_X0Y7_B_I));

wire Tile_X10Y7_RAM2FAB_D0_O0, Tile_X10Y7_RAM2FAB_D0_O1, Tile_X10Y7_RAM2FAB_D0_O2, Tile_X10Y7_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X10Y7_A (.O0(Tile_X10Y7_RAM2FAB_D0_O0), .O1(Tile_X10Y7_RAM2FAB_D0_O1), .O2(Tile_X10Y7_RAM2FAB_D0_O2), .O3(Tile_X10Y7_RAM2FAB_D0_O3));

wire Tile_X10Y7_RAM2FAB_D1_O0, Tile_X10Y7_RAM2FAB_D1_O1, Tile_X10Y7_RAM2FAB_D1_O2, Tile_X10Y7_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X10Y7_B (.O0(Tile_X10Y7_RAM2FAB_D1_O0), .O1(Tile_X10Y7_RAM2FAB_D1_O1), .O2(Tile_X10Y7_RAM2FAB_D1_O2), .O3(Tile_X10Y7_RAM2FAB_D1_O3));

wire Tile_X10Y7_RAM2FAB_D2_O0, Tile_X10Y7_RAM2FAB_D2_O1, Tile_X10Y7_RAM2FAB_D2_O2, Tile_X10Y7_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X10Y7_C (.O0(Tile_X10Y7_RAM2FAB_D2_O0), .O1(Tile_X10Y7_RAM2FAB_D2_O1), .O2(Tile_X10Y7_RAM2FAB_D2_O2), .O3(Tile_X10Y7_RAM2FAB_D2_O3));

wire Tile_X10Y7_RAM2FAB_D3_O0, Tile_X10Y7_RAM2FAB_D3_O1, Tile_X10Y7_RAM2FAB_D3_O2, Tile_X10Y7_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X10Y7_D (.O0(Tile_X10Y7_RAM2FAB_D3_O0), .O1(Tile_X10Y7_RAM2FAB_D3_O1), .O2(Tile_X10Y7_RAM2FAB_D3_O2), .O3(Tile_X10Y7_RAM2FAB_D3_O3));

wire Tile_X10Y7_FAB2RAM_D0_I0, Tile_X10Y7_FAB2RAM_D0_I1, Tile_X10Y7_FAB2RAM_D0_I2, Tile_X10Y7_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y7_E (.I0(Tile_X10Y7_FAB2RAM_D0_I0), .I1(Tile_X10Y7_FAB2RAM_D0_I1), .I2(Tile_X10Y7_FAB2RAM_D0_I2), .I3(Tile_X10Y7_FAB2RAM_D0_I3));

wire Tile_X10Y7_FAB2RAM_D1_I0, Tile_X10Y7_FAB2RAM_D1_I1, Tile_X10Y7_FAB2RAM_D1_I2, Tile_X10Y7_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y7_F (.I0(Tile_X10Y7_FAB2RAM_D1_I0), .I1(Tile_X10Y7_FAB2RAM_D1_I1), .I2(Tile_X10Y7_FAB2RAM_D1_I2), .I3(Tile_X10Y7_FAB2RAM_D1_I3));

wire Tile_X10Y7_FAB2RAM_D2_I0, Tile_X10Y7_FAB2RAM_D2_I1, Tile_X10Y7_FAB2RAM_D2_I2, Tile_X10Y7_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X10Y7_G (.I0(Tile_X10Y7_FAB2RAM_D2_I0), .I1(Tile_X10Y7_FAB2RAM_D2_I1), .I2(Tile_X10Y7_FAB2RAM_D2_I2), .I3(Tile_X10Y7_FAB2RAM_D2_I3));

wire Tile_X10Y7_FAB2RAM_D3_I0, Tile_X10Y7_FAB2RAM_D3_I1, Tile_X10Y7_FAB2RAM_D3_I2, Tile_X10Y7_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X10Y7_H (.I0(Tile_X10Y7_FAB2RAM_D3_I0), .I1(Tile_X10Y7_FAB2RAM_D3_I1), .I2(Tile_X10Y7_FAB2RAM_D3_I2), .I3(Tile_X10Y7_FAB2RAM_D3_I3));

wire Tile_X10Y7_FAB2RAM_A0_I0, Tile_X10Y7_FAB2RAM_A0_I1, Tile_X10Y7_FAB2RAM_A0_I2, Tile_X10Y7_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y7_I (.I0(Tile_X10Y7_FAB2RAM_A0_I0), .I1(Tile_X10Y7_FAB2RAM_A0_I1), .I2(Tile_X10Y7_FAB2RAM_A0_I2), .I3(Tile_X10Y7_FAB2RAM_A0_I3));

wire Tile_X10Y7_FAB2RAM_A1_I0, Tile_X10Y7_FAB2RAM_A1_I1, Tile_X10Y7_FAB2RAM_A1_I2, Tile_X10Y7_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y7_J (.I0(Tile_X10Y7_FAB2RAM_A1_I0), .I1(Tile_X10Y7_FAB2RAM_A1_I1), .I2(Tile_X10Y7_FAB2RAM_A1_I2), .I3(Tile_X10Y7_FAB2RAM_A1_I3));

wire Tile_X10Y7_FAB2RAM_C_I0, Tile_X10Y7_FAB2RAM_C_I1, Tile_X10Y7_FAB2RAM_C_I2, Tile_X10Y7_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X10Y7_K (.I0(Tile_X10Y7_FAB2RAM_C_I0), .I1(Tile_X10Y7_FAB2RAM_C_I1), .I2(Tile_X10Y7_FAB2RAM_C_I2), .I3(Tile_X10Y7_FAB2RAM_C_I3));

wire Tile_X0Y8_A_I, Tile_X0Y8_A_T, Tile_X0Y8_A_O, Tile_X0Y8_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y8_A (.O(Tile_X0Y8_A_O), .Q(Tile_X0Y8_A_Q), .I(Tile_X0Y8_A_I));

wire Tile_X0Y8_B_I, Tile_X0Y8_B_T, Tile_X0Y8_B_O, Tile_X0Y8_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y8_B (.O(Tile_X0Y8_B_O), .Q(Tile_X0Y8_B_Q), .I(Tile_X0Y8_B_I));

wire Tile_X10Y8_RAM2FAB_D0_O0, Tile_X10Y8_RAM2FAB_D0_O1, Tile_X10Y8_RAM2FAB_D0_O2, Tile_X10Y8_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X10Y8_A (.O0(Tile_X10Y8_RAM2FAB_D0_O0), .O1(Tile_X10Y8_RAM2FAB_D0_O1), .O2(Tile_X10Y8_RAM2FAB_D0_O2), .O3(Tile_X10Y8_RAM2FAB_D0_O3));

wire Tile_X10Y8_RAM2FAB_D1_O0, Tile_X10Y8_RAM2FAB_D1_O1, Tile_X10Y8_RAM2FAB_D1_O2, Tile_X10Y8_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X10Y8_B (.O0(Tile_X10Y8_RAM2FAB_D1_O0), .O1(Tile_X10Y8_RAM2FAB_D1_O1), .O2(Tile_X10Y8_RAM2FAB_D1_O2), .O3(Tile_X10Y8_RAM2FAB_D1_O3));

wire Tile_X10Y8_RAM2FAB_D2_O0, Tile_X10Y8_RAM2FAB_D2_O1, Tile_X10Y8_RAM2FAB_D2_O2, Tile_X10Y8_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X10Y8_C (.O0(Tile_X10Y8_RAM2FAB_D2_O0), .O1(Tile_X10Y8_RAM2FAB_D2_O1), .O2(Tile_X10Y8_RAM2FAB_D2_O2), .O3(Tile_X10Y8_RAM2FAB_D2_O3));

wire Tile_X10Y8_RAM2FAB_D3_O0, Tile_X10Y8_RAM2FAB_D3_O1, Tile_X10Y8_RAM2FAB_D3_O2, Tile_X10Y8_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X10Y8_D (.O0(Tile_X10Y8_RAM2FAB_D3_O0), .O1(Tile_X10Y8_RAM2FAB_D3_O1), .O2(Tile_X10Y8_RAM2FAB_D3_O2), .O3(Tile_X10Y8_RAM2FAB_D3_O3));

wire Tile_X10Y8_FAB2RAM_D0_I0, Tile_X10Y8_FAB2RAM_D0_I1, Tile_X10Y8_FAB2RAM_D0_I2, Tile_X10Y8_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y8_E (.I0(Tile_X10Y8_FAB2RAM_D0_I0), .I1(Tile_X10Y8_FAB2RAM_D0_I1), .I2(Tile_X10Y8_FAB2RAM_D0_I2), .I3(Tile_X10Y8_FAB2RAM_D0_I3));

wire Tile_X10Y8_FAB2RAM_D1_I0, Tile_X10Y8_FAB2RAM_D1_I1, Tile_X10Y8_FAB2RAM_D1_I2, Tile_X10Y8_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y8_F (.I0(Tile_X10Y8_FAB2RAM_D1_I0), .I1(Tile_X10Y8_FAB2RAM_D1_I1), .I2(Tile_X10Y8_FAB2RAM_D1_I2), .I3(Tile_X10Y8_FAB2RAM_D1_I3));

wire Tile_X10Y8_FAB2RAM_D2_I0, Tile_X10Y8_FAB2RAM_D2_I1, Tile_X10Y8_FAB2RAM_D2_I2, Tile_X10Y8_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X10Y8_G (.I0(Tile_X10Y8_FAB2RAM_D2_I0), .I1(Tile_X10Y8_FAB2RAM_D2_I1), .I2(Tile_X10Y8_FAB2RAM_D2_I2), .I3(Tile_X10Y8_FAB2RAM_D2_I3));

wire Tile_X10Y8_FAB2RAM_D3_I0, Tile_X10Y8_FAB2RAM_D3_I1, Tile_X10Y8_FAB2RAM_D3_I2, Tile_X10Y8_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X10Y8_H (.I0(Tile_X10Y8_FAB2RAM_D3_I0), .I1(Tile_X10Y8_FAB2RAM_D3_I1), .I2(Tile_X10Y8_FAB2RAM_D3_I2), .I3(Tile_X10Y8_FAB2RAM_D3_I3));

wire Tile_X10Y8_FAB2RAM_A0_I0, Tile_X10Y8_FAB2RAM_A0_I1, Tile_X10Y8_FAB2RAM_A0_I2, Tile_X10Y8_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y8_I (.I0(Tile_X10Y8_FAB2RAM_A0_I0), .I1(Tile_X10Y8_FAB2RAM_A0_I1), .I2(Tile_X10Y8_FAB2RAM_A0_I2), .I3(Tile_X10Y8_FAB2RAM_A0_I3));

wire Tile_X10Y8_FAB2RAM_A1_I0, Tile_X10Y8_FAB2RAM_A1_I1, Tile_X10Y8_FAB2RAM_A1_I2, Tile_X10Y8_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y8_J (.I0(Tile_X10Y8_FAB2RAM_A1_I0), .I1(Tile_X10Y8_FAB2RAM_A1_I1), .I2(Tile_X10Y8_FAB2RAM_A1_I2), .I3(Tile_X10Y8_FAB2RAM_A1_I3));

wire Tile_X10Y8_FAB2RAM_C_I0, Tile_X10Y8_FAB2RAM_C_I1, Tile_X10Y8_FAB2RAM_C_I2, Tile_X10Y8_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X10Y8_K (.I0(Tile_X10Y8_FAB2RAM_C_I0), .I1(Tile_X10Y8_FAB2RAM_C_I1), .I2(Tile_X10Y8_FAB2RAM_C_I2), .I3(Tile_X10Y8_FAB2RAM_C_I3));

wire Tile_X0Y9_A_I, Tile_X0Y9_A_T, Tile_X0Y9_A_O, Tile_X0Y9_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y9_A (.O(Tile_X0Y9_A_O), .Q(Tile_X0Y9_A_Q), .I(Tile_X0Y9_A_I));

wire Tile_X0Y9_B_I, Tile_X0Y9_B_T, Tile_X0Y9_B_O, Tile_X0Y9_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y9_B (.O(Tile_X0Y9_B_O), .Q(Tile_X0Y9_B_Q), .I(Tile_X0Y9_B_I));

wire Tile_X10Y9_RAM2FAB_D0_O0, Tile_X10Y9_RAM2FAB_D0_O1, Tile_X10Y9_RAM2FAB_D0_O2, Tile_X10Y9_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X10Y9_A (.O0(Tile_X10Y9_RAM2FAB_D0_O0), .O1(Tile_X10Y9_RAM2FAB_D0_O1), .O2(Tile_X10Y9_RAM2FAB_D0_O2), .O3(Tile_X10Y9_RAM2FAB_D0_O3));

wire Tile_X10Y9_RAM2FAB_D1_O0, Tile_X10Y9_RAM2FAB_D1_O1, Tile_X10Y9_RAM2FAB_D1_O2, Tile_X10Y9_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X10Y9_B (.O0(Tile_X10Y9_RAM2FAB_D1_O0), .O1(Tile_X10Y9_RAM2FAB_D1_O1), .O2(Tile_X10Y9_RAM2FAB_D1_O2), .O3(Tile_X10Y9_RAM2FAB_D1_O3));

wire Tile_X10Y9_RAM2FAB_D2_O0, Tile_X10Y9_RAM2FAB_D2_O1, Tile_X10Y9_RAM2FAB_D2_O2, Tile_X10Y9_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X10Y9_C (.O0(Tile_X10Y9_RAM2FAB_D2_O0), .O1(Tile_X10Y9_RAM2FAB_D2_O1), .O2(Tile_X10Y9_RAM2FAB_D2_O2), .O3(Tile_X10Y9_RAM2FAB_D2_O3));

wire Tile_X10Y9_RAM2FAB_D3_O0, Tile_X10Y9_RAM2FAB_D3_O1, Tile_X10Y9_RAM2FAB_D3_O2, Tile_X10Y9_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X10Y9_D (.O0(Tile_X10Y9_RAM2FAB_D3_O0), .O1(Tile_X10Y9_RAM2FAB_D3_O1), .O2(Tile_X10Y9_RAM2FAB_D3_O2), .O3(Tile_X10Y9_RAM2FAB_D3_O3));

wire Tile_X10Y9_FAB2RAM_D0_I0, Tile_X10Y9_FAB2RAM_D0_I1, Tile_X10Y9_FAB2RAM_D0_I2, Tile_X10Y9_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y9_E (.I0(Tile_X10Y9_FAB2RAM_D0_I0), .I1(Tile_X10Y9_FAB2RAM_D0_I1), .I2(Tile_X10Y9_FAB2RAM_D0_I2), .I3(Tile_X10Y9_FAB2RAM_D0_I3));

wire Tile_X10Y9_FAB2RAM_D1_I0, Tile_X10Y9_FAB2RAM_D1_I1, Tile_X10Y9_FAB2RAM_D1_I2, Tile_X10Y9_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y9_F (.I0(Tile_X10Y9_FAB2RAM_D1_I0), .I1(Tile_X10Y9_FAB2RAM_D1_I1), .I2(Tile_X10Y9_FAB2RAM_D1_I2), .I3(Tile_X10Y9_FAB2RAM_D1_I3));

wire Tile_X10Y9_FAB2RAM_D2_I0, Tile_X10Y9_FAB2RAM_D2_I1, Tile_X10Y9_FAB2RAM_D2_I2, Tile_X10Y9_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X10Y9_G (.I0(Tile_X10Y9_FAB2RAM_D2_I0), .I1(Tile_X10Y9_FAB2RAM_D2_I1), .I2(Tile_X10Y9_FAB2RAM_D2_I2), .I3(Tile_X10Y9_FAB2RAM_D2_I3));

wire Tile_X10Y9_FAB2RAM_D3_I0, Tile_X10Y9_FAB2RAM_D3_I1, Tile_X10Y9_FAB2RAM_D3_I2, Tile_X10Y9_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X10Y9_H (.I0(Tile_X10Y9_FAB2RAM_D3_I0), .I1(Tile_X10Y9_FAB2RAM_D3_I1), .I2(Tile_X10Y9_FAB2RAM_D3_I2), .I3(Tile_X10Y9_FAB2RAM_D3_I3));

wire Tile_X10Y9_FAB2RAM_A0_I0, Tile_X10Y9_FAB2RAM_A0_I1, Tile_X10Y9_FAB2RAM_A0_I2, Tile_X10Y9_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y9_I (.I0(Tile_X10Y9_FAB2RAM_A0_I0), .I1(Tile_X10Y9_FAB2RAM_A0_I1), .I2(Tile_X10Y9_FAB2RAM_A0_I2), .I3(Tile_X10Y9_FAB2RAM_A0_I3));

wire Tile_X10Y9_FAB2RAM_A1_I0, Tile_X10Y9_FAB2RAM_A1_I1, Tile_X10Y9_FAB2RAM_A1_I2, Tile_X10Y9_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y9_J (.I0(Tile_X10Y9_FAB2RAM_A1_I0), .I1(Tile_X10Y9_FAB2RAM_A1_I1), .I2(Tile_X10Y9_FAB2RAM_A1_I2), .I3(Tile_X10Y9_FAB2RAM_A1_I3));

wire Tile_X10Y9_FAB2RAM_C_I0, Tile_X10Y9_FAB2RAM_C_I1, Tile_X10Y9_FAB2RAM_C_I2, Tile_X10Y9_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X10Y9_K (.I0(Tile_X10Y9_FAB2RAM_C_I0), .I1(Tile_X10Y9_FAB2RAM_C_I1), .I2(Tile_X10Y9_FAB2RAM_C_I2), .I3(Tile_X10Y9_FAB2RAM_C_I3));

wire Tile_X0Y10_A_I, Tile_X0Y10_A_T, Tile_X0Y10_A_O, Tile_X0Y10_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y10_A (.O(Tile_X0Y10_A_O), .Q(Tile_X0Y10_A_Q), .I(Tile_X0Y10_A_I));

wire Tile_X0Y10_B_I, Tile_X0Y10_B_T, Tile_X0Y10_B_O, Tile_X0Y10_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y10_B (.O(Tile_X0Y10_B_O), .Q(Tile_X0Y10_B_Q), .I(Tile_X0Y10_B_I));

wire Tile_X10Y10_RAM2FAB_D0_O0, Tile_X10Y10_RAM2FAB_D0_O1, Tile_X10Y10_RAM2FAB_D0_O2, Tile_X10Y10_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X10Y10_A (.O0(Tile_X10Y10_RAM2FAB_D0_O0), .O1(Tile_X10Y10_RAM2FAB_D0_O1), .O2(Tile_X10Y10_RAM2FAB_D0_O2), .O3(Tile_X10Y10_RAM2FAB_D0_O3));

wire Tile_X10Y10_RAM2FAB_D1_O0, Tile_X10Y10_RAM2FAB_D1_O1, Tile_X10Y10_RAM2FAB_D1_O2, Tile_X10Y10_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X10Y10_B (.O0(Tile_X10Y10_RAM2FAB_D1_O0), .O1(Tile_X10Y10_RAM2FAB_D1_O1), .O2(Tile_X10Y10_RAM2FAB_D1_O2), .O3(Tile_X10Y10_RAM2FAB_D1_O3));

wire Tile_X10Y10_RAM2FAB_D2_O0, Tile_X10Y10_RAM2FAB_D2_O1, Tile_X10Y10_RAM2FAB_D2_O2, Tile_X10Y10_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X10Y10_C (.O0(Tile_X10Y10_RAM2FAB_D2_O0), .O1(Tile_X10Y10_RAM2FAB_D2_O1), .O2(Tile_X10Y10_RAM2FAB_D2_O2), .O3(Tile_X10Y10_RAM2FAB_D2_O3));

wire Tile_X10Y10_RAM2FAB_D3_O0, Tile_X10Y10_RAM2FAB_D3_O1, Tile_X10Y10_RAM2FAB_D3_O2, Tile_X10Y10_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X10Y10_D (.O0(Tile_X10Y10_RAM2FAB_D3_O0), .O1(Tile_X10Y10_RAM2FAB_D3_O1), .O2(Tile_X10Y10_RAM2FAB_D3_O2), .O3(Tile_X10Y10_RAM2FAB_D3_O3));

wire Tile_X10Y10_FAB2RAM_D0_I0, Tile_X10Y10_FAB2RAM_D0_I1, Tile_X10Y10_FAB2RAM_D0_I2, Tile_X10Y10_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y10_E (.I0(Tile_X10Y10_FAB2RAM_D0_I0), .I1(Tile_X10Y10_FAB2RAM_D0_I1), .I2(Tile_X10Y10_FAB2RAM_D0_I2), .I3(Tile_X10Y10_FAB2RAM_D0_I3));

wire Tile_X10Y10_FAB2RAM_D1_I0, Tile_X10Y10_FAB2RAM_D1_I1, Tile_X10Y10_FAB2RAM_D1_I2, Tile_X10Y10_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y10_F (.I0(Tile_X10Y10_FAB2RAM_D1_I0), .I1(Tile_X10Y10_FAB2RAM_D1_I1), .I2(Tile_X10Y10_FAB2RAM_D1_I2), .I3(Tile_X10Y10_FAB2RAM_D1_I3));

wire Tile_X10Y10_FAB2RAM_D2_I0, Tile_X10Y10_FAB2RAM_D2_I1, Tile_X10Y10_FAB2RAM_D2_I2, Tile_X10Y10_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X10Y10_G (.I0(Tile_X10Y10_FAB2RAM_D2_I0), .I1(Tile_X10Y10_FAB2RAM_D2_I1), .I2(Tile_X10Y10_FAB2RAM_D2_I2), .I3(Tile_X10Y10_FAB2RAM_D2_I3));

wire Tile_X10Y10_FAB2RAM_D3_I0, Tile_X10Y10_FAB2RAM_D3_I1, Tile_X10Y10_FAB2RAM_D3_I2, Tile_X10Y10_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X10Y10_H (.I0(Tile_X10Y10_FAB2RAM_D3_I0), .I1(Tile_X10Y10_FAB2RAM_D3_I1), .I2(Tile_X10Y10_FAB2RAM_D3_I2), .I3(Tile_X10Y10_FAB2RAM_D3_I3));

wire Tile_X10Y10_FAB2RAM_A0_I0, Tile_X10Y10_FAB2RAM_A0_I1, Tile_X10Y10_FAB2RAM_A0_I2, Tile_X10Y10_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y10_I (.I0(Tile_X10Y10_FAB2RAM_A0_I0), .I1(Tile_X10Y10_FAB2RAM_A0_I1), .I2(Tile_X10Y10_FAB2RAM_A0_I2), .I3(Tile_X10Y10_FAB2RAM_A0_I3));

wire Tile_X10Y10_FAB2RAM_A1_I0, Tile_X10Y10_FAB2RAM_A1_I1, Tile_X10Y10_FAB2RAM_A1_I2, Tile_X10Y10_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y10_J (.I0(Tile_X10Y10_FAB2RAM_A1_I0), .I1(Tile_X10Y10_FAB2RAM_A1_I1), .I2(Tile_X10Y10_FAB2RAM_A1_I2), .I3(Tile_X10Y10_FAB2RAM_A1_I3));

wire Tile_X10Y10_FAB2RAM_C_I0, Tile_X10Y10_FAB2RAM_C_I1, Tile_X10Y10_FAB2RAM_C_I2, Tile_X10Y10_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X10Y10_K (.I0(Tile_X10Y10_FAB2RAM_C_I0), .I1(Tile_X10Y10_FAB2RAM_C_I1), .I2(Tile_X10Y10_FAB2RAM_C_I2), .I3(Tile_X10Y10_FAB2RAM_C_I3));

wire Tile_X0Y11_A_I, Tile_X0Y11_A_T, Tile_X0Y11_A_O, Tile_X0Y11_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y11_A (.O(Tile_X0Y11_A_O), .Q(Tile_X0Y11_A_Q), .I(Tile_X0Y11_A_I));

wire Tile_X0Y11_B_I, Tile_X0Y11_B_T, Tile_X0Y11_B_O, Tile_X0Y11_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y11_B (.O(Tile_X0Y11_B_O), .Q(Tile_X0Y11_B_Q), .I(Tile_X0Y11_B_I));

wire Tile_X10Y11_RAM2FAB_D0_O0, Tile_X10Y11_RAM2FAB_D0_O1, Tile_X10Y11_RAM2FAB_D0_O2, Tile_X10Y11_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X10Y11_A (.O0(Tile_X10Y11_RAM2FAB_D0_O0), .O1(Tile_X10Y11_RAM2FAB_D0_O1), .O2(Tile_X10Y11_RAM2FAB_D0_O2), .O3(Tile_X10Y11_RAM2FAB_D0_O3));

wire Tile_X10Y11_RAM2FAB_D1_O0, Tile_X10Y11_RAM2FAB_D1_O1, Tile_X10Y11_RAM2FAB_D1_O2, Tile_X10Y11_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X10Y11_B (.O0(Tile_X10Y11_RAM2FAB_D1_O0), .O1(Tile_X10Y11_RAM2FAB_D1_O1), .O2(Tile_X10Y11_RAM2FAB_D1_O2), .O3(Tile_X10Y11_RAM2FAB_D1_O3));

wire Tile_X10Y11_RAM2FAB_D2_O0, Tile_X10Y11_RAM2FAB_D2_O1, Tile_X10Y11_RAM2FAB_D2_O2, Tile_X10Y11_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X10Y11_C (.O0(Tile_X10Y11_RAM2FAB_D2_O0), .O1(Tile_X10Y11_RAM2FAB_D2_O1), .O2(Tile_X10Y11_RAM2FAB_D2_O2), .O3(Tile_X10Y11_RAM2FAB_D2_O3));

wire Tile_X10Y11_RAM2FAB_D3_O0, Tile_X10Y11_RAM2FAB_D3_O1, Tile_X10Y11_RAM2FAB_D3_O2, Tile_X10Y11_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X10Y11_D (.O0(Tile_X10Y11_RAM2FAB_D3_O0), .O1(Tile_X10Y11_RAM2FAB_D3_O1), .O2(Tile_X10Y11_RAM2FAB_D3_O2), .O3(Tile_X10Y11_RAM2FAB_D3_O3));

wire Tile_X10Y11_FAB2RAM_D0_I0, Tile_X10Y11_FAB2RAM_D0_I1, Tile_X10Y11_FAB2RAM_D0_I2, Tile_X10Y11_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y11_E (.I0(Tile_X10Y11_FAB2RAM_D0_I0), .I1(Tile_X10Y11_FAB2RAM_D0_I1), .I2(Tile_X10Y11_FAB2RAM_D0_I2), .I3(Tile_X10Y11_FAB2RAM_D0_I3));

wire Tile_X10Y11_FAB2RAM_D1_I0, Tile_X10Y11_FAB2RAM_D1_I1, Tile_X10Y11_FAB2RAM_D1_I2, Tile_X10Y11_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y11_F (.I0(Tile_X10Y11_FAB2RAM_D1_I0), .I1(Tile_X10Y11_FAB2RAM_D1_I1), .I2(Tile_X10Y11_FAB2RAM_D1_I2), .I3(Tile_X10Y11_FAB2RAM_D1_I3));

wire Tile_X10Y11_FAB2RAM_D2_I0, Tile_X10Y11_FAB2RAM_D2_I1, Tile_X10Y11_FAB2RAM_D2_I2, Tile_X10Y11_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X10Y11_G (.I0(Tile_X10Y11_FAB2RAM_D2_I0), .I1(Tile_X10Y11_FAB2RAM_D2_I1), .I2(Tile_X10Y11_FAB2RAM_D2_I2), .I3(Tile_X10Y11_FAB2RAM_D2_I3));

wire Tile_X10Y11_FAB2RAM_D3_I0, Tile_X10Y11_FAB2RAM_D3_I1, Tile_X10Y11_FAB2RAM_D3_I2, Tile_X10Y11_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X10Y11_H (.I0(Tile_X10Y11_FAB2RAM_D3_I0), .I1(Tile_X10Y11_FAB2RAM_D3_I1), .I2(Tile_X10Y11_FAB2RAM_D3_I2), .I3(Tile_X10Y11_FAB2RAM_D3_I3));

wire Tile_X10Y11_FAB2RAM_A0_I0, Tile_X10Y11_FAB2RAM_A0_I1, Tile_X10Y11_FAB2RAM_A0_I2, Tile_X10Y11_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y11_I (.I0(Tile_X10Y11_FAB2RAM_A0_I0), .I1(Tile_X10Y11_FAB2RAM_A0_I1), .I2(Tile_X10Y11_FAB2RAM_A0_I2), .I3(Tile_X10Y11_FAB2RAM_A0_I3));

wire Tile_X10Y11_FAB2RAM_A1_I0, Tile_X10Y11_FAB2RAM_A1_I1, Tile_X10Y11_FAB2RAM_A1_I2, Tile_X10Y11_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y11_J (.I0(Tile_X10Y11_FAB2RAM_A1_I0), .I1(Tile_X10Y11_FAB2RAM_A1_I1), .I2(Tile_X10Y11_FAB2RAM_A1_I2), .I3(Tile_X10Y11_FAB2RAM_A1_I3));

wire Tile_X10Y11_FAB2RAM_C_I0, Tile_X10Y11_FAB2RAM_C_I1, Tile_X10Y11_FAB2RAM_C_I2, Tile_X10Y11_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X10Y11_K (.I0(Tile_X10Y11_FAB2RAM_C_I0), .I1(Tile_X10Y11_FAB2RAM_C_I1), .I2(Tile_X10Y11_FAB2RAM_C_I2), .I3(Tile_X10Y11_FAB2RAM_C_I3));

wire Tile_X0Y12_A_I, Tile_X0Y12_A_T, Tile_X0Y12_A_O, Tile_X0Y12_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y12_A (.O(Tile_X0Y12_A_O), .Q(Tile_X0Y12_A_Q), .I(Tile_X0Y12_A_I));

wire Tile_X0Y12_B_I, Tile_X0Y12_B_T, Tile_X0Y12_B_O, Tile_X0Y12_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y12_B (.O(Tile_X0Y12_B_O), .Q(Tile_X0Y12_B_Q), .I(Tile_X0Y12_B_I));

wire Tile_X10Y12_RAM2FAB_D0_O0, Tile_X10Y12_RAM2FAB_D0_O1, Tile_X10Y12_RAM2FAB_D0_O2, Tile_X10Y12_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X10Y12_A (.O0(Tile_X10Y12_RAM2FAB_D0_O0), .O1(Tile_X10Y12_RAM2FAB_D0_O1), .O2(Tile_X10Y12_RAM2FAB_D0_O2), .O3(Tile_X10Y12_RAM2FAB_D0_O3));

wire Tile_X10Y12_RAM2FAB_D1_O0, Tile_X10Y12_RAM2FAB_D1_O1, Tile_X10Y12_RAM2FAB_D1_O2, Tile_X10Y12_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X10Y12_B (.O0(Tile_X10Y12_RAM2FAB_D1_O0), .O1(Tile_X10Y12_RAM2FAB_D1_O1), .O2(Tile_X10Y12_RAM2FAB_D1_O2), .O3(Tile_X10Y12_RAM2FAB_D1_O3));

wire Tile_X10Y12_RAM2FAB_D2_O0, Tile_X10Y12_RAM2FAB_D2_O1, Tile_X10Y12_RAM2FAB_D2_O2, Tile_X10Y12_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X10Y12_C (.O0(Tile_X10Y12_RAM2FAB_D2_O0), .O1(Tile_X10Y12_RAM2FAB_D2_O1), .O2(Tile_X10Y12_RAM2FAB_D2_O2), .O3(Tile_X10Y12_RAM2FAB_D2_O3));

wire Tile_X10Y12_RAM2FAB_D3_O0, Tile_X10Y12_RAM2FAB_D3_O1, Tile_X10Y12_RAM2FAB_D3_O2, Tile_X10Y12_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X10Y12_D (.O0(Tile_X10Y12_RAM2FAB_D3_O0), .O1(Tile_X10Y12_RAM2FAB_D3_O1), .O2(Tile_X10Y12_RAM2FAB_D3_O2), .O3(Tile_X10Y12_RAM2FAB_D3_O3));

wire Tile_X10Y12_FAB2RAM_D0_I0, Tile_X10Y12_FAB2RAM_D0_I1, Tile_X10Y12_FAB2RAM_D0_I2, Tile_X10Y12_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y12_E (.I0(Tile_X10Y12_FAB2RAM_D0_I0), .I1(Tile_X10Y12_FAB2RAM_D0_I1), .I2(Tile_X10Y12_FAB2RAM_D0_I2), .I3(Tile_X10Y12_FAB2RAM_D0_I3));

wire Tile_X10Y12_FAB2RAM_D1_I0, Tile_X10Y12_FAB2RAM_D1_I1, Tile_X10Y12_FAB2RAM_D1_I2, Tile_X10Y12_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y12_F (.I0(Tile_X10Y12_FAB2RAM_D1_I0), .I1(Tile_X10Y12_FAB2RAM_D1_I1), .I2(Tile_X10Y12_FAB2RAM_D1_I2), .I3(Tile_X10Y12_FAB2RAM_D1_I3));

wire Tile_X10Y12_FAB2RAM_D2_I0, Tile_X10Y12_FAB2RAM_D2_I1, Tile_X10Y12_FAB2RAM_D2_I2, Tile_X10Y12_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X10Y12_G (.I0(Tile_X10Y12_FAB2RAM_D2_I0), .I1(Tile_X10Y12_FAB2RAM_D2_I1), .I2(Tile_X10Y12_FAB2RAM_D2_I2), .I3(Tile_X10Y12_FAB2RAM_D2_I3));

wire Tile_X10Y12_FAB2RAM_D3_I0, Tile_X10Y12_FAB2RAM_D3_I1, Tile_X10Y12_FAB2RAM_D3_I2, Tile_X10Y12_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X10Y12_H (.I0(Tile_X10Y12_FAB2RAM_D3_I0), .I1(Tile_X10Y12_FAB2RAM_D3_I1), .I2(Tile_X10Y12_FAB2RAM_D3_I2), .I3(Tile_X10Y12_FAB2RAM_D3_I3));

wire Tile_X10Y12_FAB2RAM_A0_I0, Tile_X10Y12_FAB2RAM_A0_I1, Tile_X10Y12_FAB2RAM_A0_I2, Tile_X10Y12_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y12_I (.I0(Tile_X10Y12_FAB2RAM_A0_I0), .I1(Tile_X10Y12_FAB2RAM_A0_I1), .I2(Tile_X10Y12_FAB2RAM_A0_I2), .I3(Tile_X10Y12_FAB2RAM_A0_I3));

wire Tile_X10Y12_FAB2RAM_A1_I0, Tile_X10Y12_FAB2RAM_A1_I1, Tile_X10Y12_FAB2RAM_A1_I2, Tile_X10Y12_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y12_J (.I0(Tile_X10Y12_FAB2RAM_A1_I0), .I1(Tile_X10Y12_FAB2RAM_A1_I1), .I2(Tile_X10Y12_FAB2RAM_A1_I2), .I3(Tile_X10Y12_FAB2RAM_A1_I3));

wire Tile_X10Y12_FAB2RAM_C_I0, Tile_X10Y12_FAB2RAM_C_I1, Tile_X10Y12_FAB2RAM_C_I2, Tile_X10Y12_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X10Y12_K (.I0(Tile_X10Y12_FAB2RAM_C_I0), .I1(Tile_X10Y12_FAB2RAM_C_I1), .I2(Tile_X10Y12_FAB2RAM_C_I2), .I3(Tile_X10Y12_FAB2RAM_C_I3));

wire Tile_X0Y13_A_I, Tile_X0Y13_A_T, Tile_X0Y13_A_O, Tile_X0Y13_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y13_A (.O(Tile_X0Y13_A_O), .Q(Tile_X0Y13_A_Q), .I(Tile_X0Y13_A_I));

wire Tile_X0Y13_B_I, Tile_X0Y13_B_T, Tile_X0Y13_B_O, Tile_X0Y13_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y13_B (.O(Tile_X0Y13_B_O), .Q(Tile_X0Y13_B_Q), .I(Tile_X0Y13_B_I));

wire Tile_X10Y13_RAM2FAB_D0_O0, Tile_X10Y13_RAM2FAB_D0_O1, Tile_X10Y13_RAM2FAB_D0_O2, Tile_X10Y13_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X10Y13_A (.O0(Tile_X10Y13_RAM2FAB_D0_O0), .O1(Tile_X10Y13_RAM2FAB_D0_O1), .O2(Tile_X10Y13_RAM2FAB_D0_O2), .O3(Tile_X10Y13_RAM2FAB_D0_O3));

wire Tile_X10Y13_RAM2FAB_D1_O0, Tile_X10Y13_RAM2FAB_D1_O1, Tile_X10Y13_RAM2FAB_D1_O2, Tile_X10Y13_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X10Y13_B (.O0(Tile_X10Y13_RAM2FAB_D1_O0), .O1(Tile_X10Y13_RAM2FAB_D1_O1), .O2(Tile_X10Y13_RAM2FAB_D1_O2), .O3(Tile_X10Y13_RAM2FAB_D1_O3));

wire Tile_X10Y13_RAM2FAB_D2_O0, Tile_X10Y13_RAM2FAB_D2_O1, Tile_X10Y13_RAM2FAB_D2_O2, Tile_X10Y13_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X10Y13_C (.O0(Tile_X10Y13_RAM2FAB_D2_O0), .O1(Tile_X10Y13_RAM2FAB_D2_O1), .O2(Tile_X10Y13_RAM2FAB_D2_O2), .O3(Tile_X10Y13_RAM2FAB_D2_O3));

wire Tile_X10Y13_RAM2FAB_D3_O0, Tile_X10Y13_RAM2FAB_D3_O1, Tile_X10Y13_RAM2FAB_D3_O2, Tile_X10Y13_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X10Y13_D (.O0(Tile_X10Y13_RAM2FAB_D3_O0), .O1(Tile_X10Y13_RAM2FAB_D3_O1), .O2(Tile_X10Y13_RAM2FAB_D3_O2), .O3(Tile_X10Y13_RAM2FAB_D3_O3));

wire Tile_X10Y13_FAB2RAM_D0_I0, Tile_X10Y13_FAB2RAM_D0_I1, Tile_X10Y13_FAB2RAM_D0_I2, Tile_X10Y13_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y13_E (.I0(Tile_X10Y13_FAB2RAM_D0_I0), .I1(Tile_X10Y13_FAB2RAM_D0_I1), .I2(Tile_X10Y13_FAB2RAM_D0_I2), .I3(Tile_X10Y13_FAB2RAM_D0_I3));

wire Tile_X10Y13_FAB2RAM_D1_I0, Tile_X10Y13_FAB2RAM_D1_I1, Tile_X10Y13_FAB2RAM_D1_I2, Tile_X10Y13_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y13_F (.I0(Tile_X10Y13_FAB2RAM_D1_I0), .I1(Tile_X10Y13_FAB2RAM_D1_I1), .I2(Tile_X10Y13_FAB2RAM_D1_I2), .I3(Tile_X10Y13_FAB2RAM_D1_I3));

wire Tile_X10Y13_FAB2RAM_D2_I0, Tile_X10Y13_FAB2RAM_D2_I1, Tile_X10Y13_FAB2RAM_D2_I2, Tile_X10Y13_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X10Y13_G (.I0(Tile_X10Y13_FAB2RAM_D2_I0), .I1(Tile_X10Y13_FAB2RAM_D2_I1), .I2(Tile_X10Y13_FAB2RAM_D2_I2), .I3(Tile_X10Y13_FAB2RAM_D2_I3));

wire Tile_X10Y13_FAB2RAM_D3_I0, Tile_X10Y13_FAB2RAM_D3_I1, Tile_X10Y13_FAB2RAM_D3_I2, Tile_X10Y13_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X10Y13_H (.I0(Tile_X10Y13_FAB2RAM_D3_I0), .I1(Tile_X10Y13_FAB2RAM_D3_I1), .I2(Tile_X10Y13_FAB2RAM_D3_I2), .I3(Tile_X10Y13_FAB2RAM_D3_I3));

wire Tile_X10Y13_FAB2RAM_A0_I0, Tile_X10Y13_FAB2RAM_A0_I1, Tile_X10Y13_FAB2RAM_A0_I2, Tile_X10Y13_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y13_I (.I0(Tile_X10Y13_FAB2RAM_A0_I0), .I1(Tile_X10Y13_FAB2RAM_A0_I1), .I2(Tile_X10Y13_FAB2RAM_A0_I2), .I3(Tile_X10Y13_FAB2RAM_A0_I3));

wire Tile_X10Y13_FAB2RAM_A1_I0, Tile_X10Y13_FAB2RAM_A1_I1, Tile_X10Y13_FAB2RAM_A1_I2, Tile_X10Y13_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y13_J (.I0(Tile_X10Y13_FAB2RAM_A1_I0), .I1(Tile_X10Y13_FAB2RAM_A1_I1), .I2(Tile_X10Y13_FAB2RAM_A1_I2), .I3(Tile_X10Y13_FAB2RAM_A1_I3));

wire Tile_X10Y13_FAB2RAM_C_I0, Tile_X10Y13_FAB2RAM_C_I1, Tile_X10Y13_FAB2RAM_C_I2, Tile_X10Y13_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X10Y13_K (.I0(Tile_X10Y13_FAB2RAM_C_I0), .I1(Tile_X10Y13_FAB2RAM_C_I1), .I2(Tile_X10Y13_FAB2RAM_C_I2), .I3(Tile_X10Y13_FAB2RAM_C_I3));

wire Tile_X0Y14_A_I, Tile_X0Y14_A_T, Tile_X0Y14_A_O, Tile_X0Y14_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y14_A (.O(Tile_X0Y14_A_O), .Q(Tile_X0Y14_A_Q), .I(Tile_X0Y14_A_I));

wire Tile_X0Y14_B_I, Tile_X0Y14_B_T, Tile_X0Y14_B_O, Tile_X0Y14_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y14_B (.O(Tile_X0Y14_B_O), .Q(Tile_X0Y14_B_Q), .I(Tile_X0Y14_B_I));

wire Tile_X10Y14_RAM2FAB_D0_O0, Tile_X10Y14_RAM2FAB_D0_O1, Tile_X10Y14_RAM2FAB_D0_O2, Tile_X10Y14_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X10Y14_A (.O0(Tile_X10Y14_RAM2FAB_D0_O0), .O1(Tile_X10Y14_RAM2FAB_D0_O1), .O2(Tile_X10Y14_RAM2FAB_D0_O2), .O3(Tile_X10Y14_RAM2FAB_D0_O3));

wire Tile_X10Y14_RAM2FAB_D1_O0, Tile_X10Y14_RAM2FAB_D1_O1, Tile_X10Y14_RAM2FAB_D1_O2, Tile_X10Y14_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X10Y14_B (.O0(Tile_X10Y14_RAM2FAB_D1_O0), .O1(Tile_X10Y14_RAM2FAB_D1_O1), .O2(Tile_X10Y14_RAM2FAB_D1_O2), .O3(Tile_X10Y14_RAM2FAB_D1_O3));

wire Tile_X10Y14_RAM2FAB_D2_O0, Tile_X10Y14_RAM2FAB_D2_O1, Tile_X10Y14_RAM2FAB_D2_O2, Tile_X10Y14_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X10Y14_C (.O0(Tile_X10Y14_RAM2FAB_D2_O0), .O1(Tile_X10Y14_RAM2FAB_D2_O1), .O2(Tile_X10Y14_RAM2FAB_D2_O2), .O3(Tile_X10Y14_RAM2FAB_D2_O3));

wire Tile_X10Y14_RAM2FAB_D3_O0, Tile_X10Y14_RAM2FAB_D3_O1, Tile_X10Y14_RAM2FAB_D3_O2, Tile_X10Y14_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X10Y14_D (.O0(Tile_X10Y14_RAM2FAB_D3_O0), .O1(Tile_X10Y14_RAM2FAB_D3_O1), .O2(Tile_X10Y14_RAM2FAB_D3_O2), .O3(Tile_X10Y14_RAM2FAB_D3_O3));

wire Tile_X10Y14_FAB2RAM_D0_I0, Tile_X10Y14_FAB2RAM_D0_I1, Tile_X10Y14_FAB2RAM_D0_I2, Tile_X10Y14_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y14_E (.I0(Tile_X10Y14_FAB2RAM_D0_I0), .I1(Tile_X10Y14_FAB2RAM_D0_I1), .I2(Tile_X10Y14_FAB2RAM_D0_I2), .I3(Tile_X10Y14_FAB2RAM_D0_I3));

wire Tile_X10Y14_FAB2RAM_D1_I0, Tile_X10Y14_FAB2RAM_D1_I1, Tile_X10Y14_FAB2RAM_D1_I2, Tile_X10Y14_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y14_F (.I0(Tile_X10Y14_FAB2RAM_D1_I0), .I1(Tile_X10Y14_FAB2RAM_D1_I1), .I2(Tile_X10Y14_FAB2RAM_D1_I2), .I3(Tile_X10Y14_FAB2RAM_D1_I3));

wire Tile_X10Y14_FAB2RAM_D2_I0, Tile_X10Y14_FAB2RAM_D2_I1, Tile_X10Y14_FAB2RAM_D2_I2, Tile_X10Y14_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X10Y14_G (.I0(Tile_X10Y14_FAB2RAM_D2_I0), .I1(Tile_X10Y14_FAB2RAM_D2_I1), .I2(Tile_X10Y14_FAB2RAM_D2_I2), .I3(Tile_X10Y14_FAB2RAM_D2_I3));

wire Tile_X10Y14_FAB2RAM_D3_I0, Tile_X10Y14_FAB2RAM_D3_I1, Tile_X10Y14_FAB2RAM_D3_I2, Tile_X10Y14_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X10Y14_H (.I0(Tile_X10Y14_FAB2RAM_D3_I0), .I1(Tile_X10Y14_FAB2RAM_D3_I1), .I2(Tile_X10Y14_FAB2RAM_D3_I2), .I3(Tile_X10Y14_FAB2RAM_D3_I3));

wire Tile_X10Y14_FAB2RAM_A0_I0, Tile_X10Y14_FAB2RAM_A0_I1, Tile_X10Y14_FAB2RAM_A0_I2, Tile_X10Y14_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y14_I (.I0(Tile_X10Y14_FAB2RAM_A0_I0), .I1(Tile_X10Y14_FAB2RAM_A0_I1), .I2(Tile_X10Y14_FAB2RAM_A0_I2), .I3(Tile_X10Y14_FAB2RAM_A0_I3));

wire Tile_X10Y14_FAB2RAM_A1_I0, Tile_X10Y14_FAB2RAM_A1_I1, Tile_X10Y14_FAB2RAM_A1_I2, Tile_X10Y14_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y14_J (.I0(Tile_X10Y14_FAB2RAM_A1_I0), .I1(Tile_X10Y14_FAB2RAM_A1_I1), .I2(Tile_X10Y14_FAB2RAM_A1_I2), .I3(Tile_X10Y14_FAB2RAM_A1_I3));

wire Tile_X10Y14_FAB2RAM_C_I0, Tile_X10Y14_FAB2RAM_C_I1, Tile_X10Y14_FAB2RAM_C_I2, Tile_X10Y14_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X10Y14_K (.I0(Tile_X10Y14_FAB2RAM_C_I0), .I1(Tile_X10Y14_FAB2RAM_C_I1), .I2(Tile_X10Y14_FAB2RAM_C_I2), .I3(Tile_X10Y14_FAB2RAM_C_I3));

wire Tile_X0Y15_A_I, Tile_X0Y15_A_T, Tile_X0Y15_A_O, Tile_X0Y15_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y15_A (.O(Tile_X0Y15_A_O), .Q(Tile_X0Y15_A_Q), .I(Tile_X0Y15_A_I));

wire Tile_X0Y15_B_I, Tile_X0Y15_B_T, Tile_X0Y15_B_O, Tile_X0Y15_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y15_B (.O(Tile_X0Y15_B_O), .Q(Tile_X0Y15_B_Q), .I(Tile_X0Y15_B_I));

wire Tile_X10Y15_RAM2FAB_D0_O0, Tile_X10Y15_RAM2FAB_D0_O1, Tile_X10Y15_RAM2FAB_D0_O2, Tile_X10Y15_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X10Y15_A (.O0(Tile_X10Y15_RAM2FAB_D0_O0), .O1(Tile_X10Y15_RAM2FAB_D0_O1), .O2(Tile_X10Y15_RAM2FAB_D0_O2), .O3(Tile_X10Y15_RAM2FAB_D0_O3));

wire Tile_X10Y15_RAM2FAB_D1_O0, Tile_X10Y15_RAM2FAB_D1_O1, Tile_X10Y15_RAM2FAB_D1_O2, Tile_X10Y15_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X10Y15_B (.O0(Tile_X10Y15_RAM2FAB_D1_O0), .O1(Tile_X10Y15_RAM2FAB_D1_O1), .O2(Tile_X10Y15_RAM2FAB_D1_O2), .O3(Tile_X10Y15_RAM2FAB_D1_O3));

wire Tile_X10Y15_RAM2FAB_D2_O0, Tile_X10Y15_RAM2FAB_D2_O1, Tile_X10Y15_RAM2FAB_D2_O2, Tile_X10Y15_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X10Y15_C (.O0(Tile_X10Y15_RAM2FAB_D2_O0), .O1(Tile_X10Y15_RAM2FAB_D2_O1), .O2(Tile_X10Y15_RAM2FAB_D2_O2), .O3(Tile_X10Y15_RAM2FAB_D2_O3));

wire Tile_X10Y15_RAM2FAB_D3_O0, Tile_X10Y15_RAM2FAB_D3_O1, Tile_X10Y15_RAM2FAB_D3_O2, Tile_X10Y15_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X10Y15_D (.O0(Tile_X10Y15_RAM2FAB_D3_O0), .O1(Tile_X10Y15_RAM2FAB_D3_O1), .O2(Tile_X10Y15_RAM2FAB_D3_O2), .O3(Tile_X10Y15_RAM2FAB_D3_O3));

wire Tile_X10Y15_FAB2RAM_D0_I0, Tile_X10Y15_FAB2RAM_D0_I1, Tile_X10Y15_FAB2RAM_D0_I2, Tile_X10Y15_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y15_E (.I0(Tile_X10Y15_FAB2RAM_D0_I0), .I1(Tile_X10Y15_FAB2RAM_D0_I1), .I2(Tile_X10Y15_FAB2RAM_D0_I2), .I3(Tile_X10Y15_FAB2RAM_D0_I3));

wire Tile_X10Y15_FAB2RAM_D1_I0, Tile_X10Y15_FAB2RAM_D1_I1, Tile_X10Y15_FAB2RAM_D1_I2, Tile_X10Y15_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y15_F (.I0(Tile_X10Y15_FAB2RAM_D1_I0), .I1(Tile_X10Y15_FAB2RAM_D1_I1), .I2(Tile_X10Y15_FAB2RAM_D1_I2), .I3(Tile_X10Y15_FAB2RAM_D1_I3));

wire Tile_X10Y15_FAB2RAM_D2_I0, Tile_X10Y15_FAB2RAM_D2_I1, Tile_X10Y15_FAB2RAM_D2_I2, Tile_X10Y15_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X10Y15_G (.I0(Tile_X10Y15_FAB2RAM_D2_I0), .I1(Tile_X10Y15_FAB2RAM_D2_I1), .I2(Tile_X10Y15_FAB2RAM_D2_I2), .I3(Tile_X10Y15_FAB2RAM_D2_I3));

wire Tile_X10Y15_FAB2RAM_D3_I0, Tile_X10Y15_FAB2RAM_D3_I1, Tile_X10Y15_FAB2RAM_D3_I2, Tile_X10Y15_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X10Y15_H (.I0(Tile_X10Y15_FAB2RAM_D3_I0), .I1(Tile_X10Y15_FAB2RAM_D3_I1), .I2(Tile_X10Y15_FAB2RAM_D3_I2), .I3(Tile_X10Y15_FAB2RAM_D3_I3));

wire Tile_X10Y15_FAB2RAM_A0_I0, Tile_X10Y15_FAB2RAM_A0_I1, Tile_X10Y15_FAB2RAM_A0_I2, Tile_X10Y15_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y15_I (.I0(Tile_X10Y15_FAB2RAM_A0_I0), .I1(Tile_X10Y15_FAB2RAM_A0_I1), .I2(Tile_X10Y15_FAB2RAM_A0_I2), .I3(Tile_X10Y15_FAB2RAM_A0_I3));

wire Tile_X10Y15_FAB2RAM_A1_I0, Tile_X10Y15_FAB2RAM_A1_I1, Tile_X10Y15_FAB2RAM_A1_I2, Tile_X10Y15_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y15_J (.I0(Tile_X10Y15_FAB2RAM_A1_I0), .I1(Tile_X10Y15_FAB2RAM_A1_I1), .I2(Tile_X10Y15_FAB2RAM_A1_I2), .I3(Tile_X10Y15_FAB2RAM_A1_I3));

wire Tile_X10Y15_FAB2RAM_C_I0, Tile_X10Y15_FAB2RAM_C_I1, Tile_X10Y15_FAB2RAM_C_I2, Tile_X10Y15_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X10Y15_K (.I0(Tile_X10Y15_FAB2RAM_C_I0), .I1(Tile_X10Y15_FAB2RAM_C_I1), .I2(Tile_X10Y15_FAB2RAM_C_I2), .I3(Tile_X10Y15_FAB2RAM_C_I3));

wire Tile_X0Y16_A_I, Tile_X0Y16_A_T, Tile_X0Y16_A_O, Tile_X0Y16_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y16_A (.O(Tile_X0Y16_A_O), .Q(Tile_X0Y16_A_Q), .I(Tile_X0Y16_A_I));

wire Tile_X0Y16_B_I, Tile_X0Y16_B_T, Tile_X0Y16_B_O, Tile_X0Y16_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y16_B (.O(Tile_X0Y16_B_O), .Q(Tile_X0Y16_B_Q), .I(Tile_X0Y16_B_I));

wire Tile_X10Y16_RAM2FAB_D0_O0, Tile_X10Y16_RAM2FAB_D0_O1, Tile_X10Y16_RAM2FAB_D0_O2, Tile_X10Y16_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X10Y16_A (.O0(Tile_X10Y16_RAM2FAB_D0_O0), .O1(Tile_X10Y16_RAM2FAB_D0_O1), .O2(Tile_X10Y16_RAM2FAB_D0_O2), .O3(Tile_X10Y16_RAM2FAB_D0_O3));

wire Tile_X10Y16_RAM2FAB_D1_O0, Tile_X10Y16_RAM2FAB_D1_O1, Tile_X10Y16_RAM2FAB_D1_O2, Tile_X10Y16_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X10Y16_B (.O0(Tile_X10Y16_RAM2FAB_D1_O0), .O1(Tile_X10Y16_RAM2FAB_D1_O1), .O2(Tile_X10Y16_RAM2FAB_D1_O2), .O3(Tile_X10Y16_RAM2FAB_D1_O3));

wire Tile_X10Y16_RAM2FAB_D2_O0, Tile_X10Y16_RAM2FAB_D2_O1, Tile_X10Y16_RAM2FAB_D2_O2, Tile_X10Y16_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X10Y16_C (.O0(Tile_X10Y16_RAM2FAB_D2_O0), .O1(Tile_X10Y16_RAM2FAB_D2_O1), .O2(Tile_X10Y16_RAM2FAB_D2_O2), .O3(Tile_X10Y16_RAM2FAB_D2_O3));

wire Tile_X10Y16_RAM2FAB_D3_O0, Tile_X10Y16_RAM2FAB_D3_O1, Tile_X10Y16_RAM2FAB_D3_O2, Tile_X10Y16_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X10Y16_D (.O0(Tile_X10Y16_RAM2FAB_D3_O0), .O1(Tile_X10Y16_RAM2FAB_D3_O1), .O2(Tile_X10Y16_RAM2FAB_D3_O2), .O3(Tile_X10Y16_RAM2FAB_D3_O3));

wire Tile_X10Y16_FAB2RAM_D0_I0, Tile_X10Y16_FAB2RAM_D0_I1, Tile_X10Y16_FAB2RAM_D0_I2, Tile_X10Y16_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y16_E (.I0(Tile_X10Y16_FAB2RAM_D0_I0), .I1(Tile_X10Y16_FAB2RAM_D0_I1), .I2(Tile_X10Y16_FAB2RAM_D0_I2), .I3(Tile_X10Y16_FAB2RAM_D0_I3));

wire Tile_X10Y16_FAB2RAM_D1_I0, Tile_X10Y16_FAB2RAM_D1_I1, Tile_X10Y16_FAB2RAM_D1_I2, Tile_X10Y16_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y16_F (.I0(Tile_X10Y16_FAB2RAM_D1_I0), .I1(Tile_X10Y16_FAB2RAM_D1_I1), .I2(Tile_X10Y16_FAB2RAM_D1_I2), .I3(Tile_X10Y16_FAB2RAM_D1_I3));

wire Tile_X10Y16_FAB2RAM_D2_I0, Tile_X10Y16_FAB2RAM_D2_I1, Tile_X10Y16_FAB2RAM_D2_I2, Tile_X10Y16_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X10Y16_G (.I0(Tile_X10Y16_FAB2RAM_D2_I0), .I1(Tile_X10Y16_FAB2RAM_D2_I1), .I2(Tile_X10Y16_FAB2RAM_D2_I2), .I3(Tile_X10Y16_FAB2RAM_D2_I3));

wire Tile_X10Y16_FAB2RAM_D3_I0, Tile_X10Y16_FAB2RAM_D3_I1, Tile_X10Y16_FAB2RAM_D3_I2, Tile_X10Y16_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X10Y16_H (.I0(Tile_X10Y16_FAB2RAM_D3_I0), .I1(Tile_X10Y16_FAB2RAM_D3_I1), .I2(Tile_X10Y16_FAB2RAM_D3_I2), .I3(Tile_X10Y16_FAB2RAM_D3_I3));

wire Tile_X10Y16_FAB2RAM_A0_I0, Tile_X10Y16_FAB2RAM_A0_I1, Tile_X10Y16_FAB2RAM_A0_I2, Tile_X10Y16_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X10Y16_I (.I0(Tile_X10Y16_FAB2RAM_A0_I0), .I1(Tile_X10Y16_FAB2RAM_A0_I1), .I2(Tile_X10Y16_FAB2RAM_A0_I2), .I3(Tile_X10Y16_FAB2RAM_A0_I3));

wire Tile_X10Y16_FAB2RAM_A1_I0, Tile_X10Y16_FAB2RAM_A1_I1, Tile_X10Y16_FAB2RAM_A1_I2, Tile_X10Y16_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X10Y16_J (.I0(Tile_X10Y16_FAB2RAM_A1_I0), .I1(Tile_X10Y16_FAB2RAM_A1_I1), .I2(Tile_X10Y16_FAB2RAM_A1_I2), .I3(Tile_X10Y16_FAB2RAM_A1_I3));

wire Tile_X10Y16_FAB2RAM_C_I0, Tile_X10Y16_FAB2RAM_C_I1, Tile_X10Y16_FAB2RAM_C_I2, Tile_X10Y16_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X10Y16_K (.I0(Tile_X10Y16_FAB2RAM_C_I0), .I1(Tile_X10Y16_FAB2RAM_C_I1), .I2(Tile_X10Y16_FAB2RAM_C_I2), .I3(Tile_X10Y16_FAB2RAM_C_I3));

endmodule