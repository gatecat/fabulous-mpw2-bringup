module eFPGA_CPU_top(wb_clk_i, wb_rst_i, wbs_stb_i, wbs_cyc_i, wbs_we_i, wbs_sel_i, wbs_dat_i, wbs_adr_i, wbs_ack_o, wbs_dat_o, la_data_out, la_data_in, io_in, io_out, io_oeb, user_clock2);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire \A_config_C[0] ;
  wire \A_config_C[10] ;
  wire \A_config_C[11] ;
  wire \A_config_C[12] ;
  wire \A_config_C[13] ;
  wire \A_config_C[14] ;
  wire \A_config_C[15] ;
  wire \A_config_C[16] ;
  wire \A_config_C[17] ;
  wire \A_config_C[18] ;
  wire \A_config_C[19] ;
  wire \A_config_C[1] ;
  wire \A_config_C[2] ;
  wire \A_config_C[3] ;
  wire \A_config_C[4] ;
  wire \A_config_C[5] ;
  wire \A_config_C[6] ;
  wire \A_config_C[7] ;
  wire \A_config_C[8] ;
  wire \A_config_C[9] ;
  wire \B_config_C[0] ;
  wire \B_config_C[10] ;
  wire \B_config_C[11] ;
  wire \B_config_C[12] ;
  wire \B_config_C[13] ;
  wire \B_config_C[14] ;
  wire \B_config_C[15] ;
  wire \B_config_C[16] ;
  wire \B_config_C[17] ;
  wire \B_config_C[18] ;
  wire \B_config_C[19] ;
  wire \B_config_C[1] ;
  wire \B_config_C[2] ;
  wire \B_config_C[3] ;
  wire \B_config_C[4] ;
  wire \B_config_C[5] ;
  wire \B_config_C[6] ;
  wire \B_config_C[7] ;
  wire \B_config_C[8] ;
  wire \B_config_C[9] ;
  wire CLK;
  wire ComActive;
  wire \Config_accessC[0] ;
  wire \Config_accessC[10] ;
  wire \Config_accessC[11] ;
  wire \Config_accessC[12] ;
  wire \Config_accessC[13] ;
  wire \Config_accessC[14] ;
  wire \Config_accessC[15] ;
  wire \Config_accessC[16] ;
  wire \Config_accessC[17] ;
  wire \Config_accessC[18] ;
  wire \Config_accessC[19] ;
  wire \Config_accessC[1] ;
  wire \Config_accessC[2] ;
  wire \Config_accessC[3] ;
  wire \Config_accessC[4] ;
  wire \Config_accessC[5] ;
  wire \Config_accessC[6] ;
  wire \Config_accessC[7] ;
  wire \Config_accessC[8] ;
  wire \Config_accessC[9] ;
  wire \E_OPA[0] ;
  wire \E_OPA[10] ;
  wire \E_OPA[11] ;
  wire \E_OPA[12] ;
  wire \E_OPA[13] ;
  wire \E_OPA[14] ;
  wire \E_OPA[15] ;
  wire \E_OPA[16] ;
  wire \E_OPA[17] ;
  wire \E_OPA[18] ;
  wire \E_OPA[19] ;
  wire \E_OPA[1] ;
  wire \E_OPA[20] ;
  wire \E_OPA[21] ;
  wire \E_OPA[22] ;
  wire \E_OPA[23] ;
  wire \E_OPA[24] ;
  wire \E_OPA[25] ;
  wire \E_OPA[26] ;
  wire \E_OPA[27] ;
  wire \E_OPA[28] ;
  wire \E_OPA[29] ;
  wire \E_OPA[2] ;
  wire \E_OPA[30] ;
  wire \E_OPA[31] ;
  wire \E_OPA[32] ;
  wire \E_OPA[33] ;
  wire \E_OPA[34] ;
  wire \E_OPA[35] ;
  wire \E_OPA[3] ;
  wire \E_OPA[4] ;
  wire \E_OPA[5] ;
  wire \E_OPA[6] ;
  wire \E_OPA[7] ;
  wire \E_OPA[8] ;
  wire \E_OPA[9] ;
  wire \E_OPB[0] ;
  wire \E_OPB[10] ;
  wire \E_OPB[11] ;
  wire \E_OPB[12] ;
  wire \E_OPB[13] ;
  wire \E_OPB[14] ;
  wire \E_OPB[15] ;
  wire \E_OPB[16] ;
  wire \E_OPB[17] ;
  wire \E_OPB[18] ;
  wire \E_OPB[19] ;
  wire \E_OPB[1] ;
  wire \E_OPB[20] ;
  wire \E_OPB[21] ;
  wire \E_OPB[22] ;
  wire \E_OPB[23] ;
  wire \E_OPB[24] ;
  wire \E_OPB[25] ;
  wire \E_OPB[26] ;
  wire \E_OPB[27] ;
  wire \E_OPB[28] ;
  wire \E_OPB[29] ;
  wire \E_OPB[2] ;
  wire \E_OPB[30] ;
  wire \E_OPB[31] ;
  wire \E_OPB[32] ;
  wire \E_OPB[33] ;
  wire \E_OPB[34] ;
  wire \E_OPB[35] ;
  wire \E_OPB[3] ;
  wire \E_OPB[4] ;
  wire \E_OPB[5] ;
  wire \E_OPB[6] ;
  wire \E_OPB[7] ;
  wire \E_OPB[8] ;
  wire \E_OPB[9] ;
  wire \E_RES0[0] ;
  wire \E_RES0[10] ;
  wire \E_RES0[11] ;
  wire \E_RES0[12] ;
  wire \E_RES0[13] ;
  wire \E_RES0[14] ;
  wire \E_RES0[15] ;
  wire \E_RES0[16] ;
  wire \E_RES0[17] ;
  wire \E_RES0[18] ;
  wire \E_RES0[19] ;
  wire \E_RES0[1] ;
  wire \E_RES0[20] ;
  wire \E_RES0[21] ;
  wire \E_RES0[22] ;
  wire \E_RES0[23] ;
  wire \E_RES0[24] ;
  wire \E_RES0[25] ;
  wire \E_RES0[26] ;
  wire \E_RES0[27] ;
  wire \E_RES0[28] ;
  wire \E_RES0[29] ;
  wire \E_RES0[2] ;
  wire \E_RES0[30] ;
  wire \E_RES0[31] ;
  wire \E_RES0[32] ;
  wire \E_RES0[33] ;
  wire \E_RES0[34] ;
  wire \E_RES0[35] ;
  wire \E_RES0[3] ;
  wire \E_RES0[4] ;
  wire \E_RES0[5] ;
  wire \E_RES0[6] ;
  wire \E_RES0[7] ;
  wire \E_RES0[8] ;
  wire \E_RES0[9] ;
  wire \E_RES1[0] ;
  wire \E_RES1[10] ;
  wire \E_RES1[11] ;
  wire \E_RES1[12] ;
  wire \E_RES1[13] ;
  wire \E_RES1[14] ;
  wire \E_RES1[15] ;
  wire \E_RES1[16] ;
  wire \E_RES1[17] ;
  wire \E_RES1[18] ;
  wire \E_RES1[19] ;
  wire \E_RES1[1] ;
  wire \E_RES1[20] ;
  wire \E_RES1[21] ;
  wire \E_RES1[22] ;
  wire \E_RES1[23] ;
  wire \E_RES1[24] ;
  wire \E_RES1[25] ;
  wire \E_RES1[26] ;
  wire \E_RES1[27] ;
  wire \E_RES1[28] ;
  wire \E_RES1[29] ;
  wire \E_RES1[2] ;
  wire \E_RES1[30] ;
  wire \E_RES1[31] ;
  wire \E_RES1[32] ;
  wire \E_RES1[33] ;
  wire \E_RES1[34] ;
  wire \E_RES1[35] ;
  wire \E_RES1[3] ;
  wire \E_RES1[4] ;
  wire \E_RES1[5] ;
  wire \E_RES1[6] ;
  wire \E_RES1[7] ;
  wire \E_RES1[8] ;
  wire \E_RES1[9] ;
  wire \E_RES2[0] ;
  wire \E_RES2[10] ;
  wire \E_RES2[11] ;
  wire \E_RES2[12] ;
  wire \E_RES2[13] ;
  wire \E_RES2[14] ;
  wire \E_RES2[15] ;
  wire \E_RES2[16] ;
  wire \E_RES2[17] ;
  wire \E_RES2[18] ;
  wire \E_RES2[19] ;
  wire \E_RES2[1] ;
  wire \E_RES2[20] ;
  wire \E_RES2[21] ;
  wire \E_RES2[22] ;
  wire \E_RES2[23] ;
  wire \E_RES2[24] ;
  wire \E_RES2[25] ;
  wire \E_RES2[26] ;
  wire \E_RES2[27] ;
  wire \E_RES2[28] ;
  wire \E_RES2[29] ;
  wire \E_RES2[2] ;
  wire \E_RES2[30] ;
  wire \E_RES2[31] ;
  wire \E_RES2[32] ;
  wire \E_RES2[33] ;
  wire \E_RES2[34] ;
  wire \E_RES2[35] ;
  wire \E_RES2[3] ;
  wire \E_RES2[4] ;
  wire \E_RES2[5] ;
  wire \E_RES2[6] ;
  wire \E_RES2[7] ;
  wire \E_RES2[8] ;
  wire \E_RES2[9] ;
  wire \FAB2RAM_A[0] ;
  wire \FAB2RAM_A[10] ;
  wire \FAB2RAM_A[11] ;
  wire \FAB2RAM_A[12] ;
  wire \FAB2RAM_A[13] ;
  wire \FAB2RAM_A[14] ;
  wire \FAB2RAM_A[15] ;
  wire \FAB2RAM_A[16] ;
  wire \FAB2RAM_A[17] ;
  wire \FAB2RAM_A[18] ;
  wire \FAB2RAM_A[19] ;
  wire \FAB2RAM_A[1] ;
  wire \FAB2RAM_A[20] ;
  wire \FAB2RAM_A[21] ;
  wire \FAB2RAM_A[22] ;
  wire \FAB2RAM_A[23] ;
  wire \FAB2RAM_A[24] ;
  wire \FAB2RAM_A[25] ;
  wire \FAB2RAM_A[26] ;
  wire \FAB2RAM_A[27] ;
  wire \FAB2RAM_A[28] ;
  wire \FAB2RAM_A[29] ;
  wire \FAB2RAM_A[2] ;
  wire \FAB2RAM_A[30] ;
  wire \FAB2RAM_A[31] ;
  wire \FAB2RAM_A[32] ;
  wire \FAB2RAM_A[33] ;
  wire \FAB2RAM_A[34] ;
  wire \FAB2RAM_A[35] ;
  wire \FAB2RAM_A[36] ;
  wire \FAB2RAM_A[37] ;
  wire \FAB2RAM_A[38] ;
  wire \FAB2RAM_A[39] ;
  wire \FAB2RAM_A[3] ;
  wire \FAB2RAM_A[4] ;
  wire \FAB2RAM_A[5] ;
  wire \FAB2RAM_A[6] ;
  wire \FAB2RAM_A[7] ;
  wire \FAB2RAM_A[8] ;
  wire \FAB2RAM_A[9] ;
  wire \FAB2RAM_C[0] ;
  wire \FAB2RAM_C[10] ;
  wire \FAB2RAM_C[11] ;
  wire \FAB2RAM_C[12] ;
  wire \FAB2RAM_C[13] ;
  wire \FAB2RAM_C[14] ;
  wire \FAB2RAM_C[15] ;
  wire \FAB2RAM_C[16] ;
  wire \FAB2RAM_C[17] ;
  wire \FAB2RAM_C[18] ;
  wire \FAB2RAM_C[19] ;
  wire \FAB2RAM_C[1] ;
  wire \FAB2RAM_C[2] ;
  wire \FAB2RAM_C[3] ;
  wire \FAB2RAM_C[4] ;
  wire \FAB2RAM_C[5] ;
  wire \FAB2RAM_C[6] ;
  wire \FAB2RAM_C[7] ;
  wire \FAB2RAM_C[8] ;
  wire \FAB2RAM_C[9] ;
  wire \FAB2RAM_D[0] ;
  wire \FAB2RAM_D[10] ;
  wire \FAB2RAM_D[11] ;
  wire \FAB2RAM_D[12] ;
  wire \FAB2RAM_D[13] ;
  wire \FAB2RAM_D[14] ;
  wire \FAB2RAM_D[15] ;
  wire \FAB2RAM_D[16] ;
  wire \FAB2RAM_D[17] ;
  wire \FAB2RAM_D[18] ;
  wire \FAB2RAM_D[19] ;
  wire \FAB2RAM_D[1] ;
  wire \FAB2RAM_D[20] ;
  wire \FAB2RAM_D[21] ;
  wire \FAB2RAM_D[22] ;
  wire \FAB2RAM_D[23] ;
  wire \FAB2RAM_D[24] ;
  wire \FAB2RAM_D[25] ;
  wire \FAB2RAM_D[26] ;
  wire \FAB2RAM_D[27] ;
  wire \FAB2RAM_D[28] ;
  wire \FAB2RAM_D[29] ;
  wire \FAB2RAM_D[2] ;
  wire \FAB2RAM_D[30] ;
  wire \FAB2RAM_D[31] ;
  wire \FAB2RAM_D[32] ;
  wire \FAB2RAM_D[33] ;
  wire \FAB2RAM_D[34] ;
  wire \FAB2RAM_D[35] ;
  wire \FAB2RAM_D[36] ;
  wire \FAB2RAM_D[37] ;
  wire \FAB2RAM_D[38] ;
  wire \FAB2RAM_D[39] ;
  wire \FAB2RAM_D[3] ;
  wire \FAB2RAM_D[40] ;
  wire \FAB2RAM_D[41] ;
  wire \FAB2RAM_D[42] ;
  wire \FAB2RAM_D[43] ;
  wire \FAB2RAM_D[44] ;
  wire \FAB2RAM_D[45] ;
  wire \FAB2RAM_D[46] ;
  wire \FAB2RAM_D[47] ;
  wire \FAB2RAM_D[48] ;
  wire \FAB2RAM_D[49] ;
  wire \FAB2RAM_D[4] ;
  wire \FAB2RAM_D[50] ;
  wire \FAB2RAM_D[51] ;
  wire \FAB2RAM_D[52] ;
  wire \FAB2RAM_D[53] ;
  wire \FAB2RAM_D[54] ;
  wire \FAB2RAM_D[55] ;
  wire \FAB2RAM_D[56] ;
  wire \FAB2RAM_D[57] ;
  wire \FAB2RAM_D[58] ;
  wire \FAB2RAM_D[59] ;
  wire \FAB2RAM_D[5] ;
  wire \FAB2RAM_D[60] ;
  wire \FAB2RAM_D[61] ;
  wire \FAB2RAM_D[62] ;
  wire \FAB2RAM_D[63] ;
  wire \FAB2RAM_D[64] ;
  wire \FAB2RAM_D[65] ;
  wire \FAB2RAM_D[66] ;
  wire \FAB2RAM_D[67] ;
  wire \FAB2RAM_D[68] ;
  wire \FAB2RAM_D[69] ;
  wire \FAB2RAM_D[6] ;
  wire \FAB2RAM_D[70] ;
  wire \FAB2RAM_D[71] ;
  wire \FAB2RAM_D[72] ;
  wire \FAB2RAM_D[73] ;
  wire \FAB2RAM_D[74] ;
  wire \FAB2RAM_D[75] ;
  wire \FAB2RAM_D[76] ;
  wire \FAB2RAM_D[77] ;
  wire \FAB2RAM_D[78] ;
  wire \FAB2RAM_D[79] ;
  wire \FAB2RAM_D[7] ;
  wire \FAB2RAM_D[8] ;
  wire \FAB2RAM_D[9] ;
  wire \FrameAddressRegister[0] ;
  wire \FrameAddressRegister[10] ;
  wire \FrameAddressRegister[11] ;
  wire \FrameAddressRegister[12] ;
  wire \FrameAddressRegister[13] ;
  wire \FrameAddressRegister[14] ;
  wire \FrameAddressRegister[15] ;
  wire \FrameAddressRegister[16] ;
  wire \FrameAddressRegister[17] ;
  wire \FrameAddressRegister[18] ;
  wire \FrameAddressRegister[19] ;
  wire \FrameAddressRegister[1] ;
  wire \FrameAddressRegister[20] ;
  wire \FrameAddressRegister[21] ;
  wire \FrameAddressRegister[22] ;
  wire \FrameAddressRegister[23] ;
  wire \FrameAddressRegister[24] ;
  wire \FrameAddressRegister[25] ;
  wire \FrameAddressRegister[26] ;
  wire \FrameAddressRegister[27] ;
  wire \FrameAddressRegister[28] ;
  wire \FrameAddressRegister[29] ;
  wire \FrameAddressRegister[2] ;
  wire \FrameAddressRegister[30] ;
  wire \FrameAddressRegister[31] ;
  wire \FrameAddressRegister[3] ;
  wire \FrameAddressRegister[4] ;
  wire \FrameAddressRegister[5] ;
  wire \FrameAddressRegister[6] ;
  wire \FrameAddressRegister[7] ;
  wire \FrameAddressRegister[8] ;
  wire \FrameAddressRegister[9] ;
  wire \FrameData[100] ;
  wire \FrameData[101] ;
  wire \FrameData[102] ;
  wire \FrameData[103] ;
  wire \FrameData[104] ;
  wire \FrameData[105] ;
  wire \FrameData[106] ;
  wire \FrameData[107] ;
  wire \FrameData[108] ;
  wire \FrameData[109] ;
  wire \FrameData[110] ;
  wire \FrameData[111] ;
  wire \FrameData[112] ;
  wire \FrameData[113] ;
  wire \FrameData[114] ;
  wire \FrameData[115] ;
  wire \FrameData[116] ;
  wire \FrameData[117] ;
  wire \FrameData[118] ;
  wire \FrameData[119] ;
  wire \FrameData[120] ;
  wire \FrameData[121] ;
  wire \FrameData[122] ;
  wire \FrameData[123] ;
  wire \FrameData[124] ;
  wire \FrameData[125] ;
  wire \FrameData[126] ;
  wire \FrameData[127] ;
  wire \FrameData[128] ;
  wire \FrameData[129] ;
  wire \FrameData[130] ;
  wire \FrameData[131] ;
  wire \FrameData[132] ;
  wire \FrameData[133] ;
  wire \FrameData[134] ;
  wire \FrameData[135] ;
  wire \FrameData[136] ;
  wire \FrameData[137] ;
  wire \FrameData[138] ;
  wire \FrameData[139] ;
  wire \FrameData[140] ;
  wire \FrameData[141] ;
  wire \FrameData[142] ;
  wire \FrameData[143] ;
  wire \FrameData[144] ;
  wire \FrameData[145] ;
  wire \FrameData[146] ;
  wire \FrameData[147] ;
  wire \FrameData[148] ;
  wire \FrameData[149] ;
  wire \FrameData[150] ;
  wire \FrameData[151] ;
  wire \FrameData[152] ;
  wire \FrameData[153] ;
  wire \FrameData[154] ;
  wire \FrameData[155] ;
  wire \FrameData[156] ;
  wire \FrameData[157] ;
  wire \FrameData[158] ;
  wire \FrameData[159] ;
  wire \FrameData[160] ;
  wire \FrameData[161] ;
  wire \FrameData[162] ;
  wire \FrameData[163] ;
  wire \FrameData[164] ;
  wire \FrameData[165] ;
  wire \FrameData[166] ;
  wire \FrameData[167] ;
  wire \FrameData[168] ;
  wire \FrameData[169] ;
  wire \FrameData[170] ;
  wire \FrameData[171] ;
  wire \FrameData[172] ;
  wire \FrameData[173] ;
  wire \FrameData[174] ;
  wire \FrameData[175] ;
  wire \FrameData[176] ;
  wire \FrameData[177] ;
  wire \FrameData[178] ;
  wire \FrameData[179] ;
  wire \FrameData[180] ;
  wire \FrameData[181] ;
  wire \FrameData[182] ;
  wire \FrameData[183] ;
  wire \FrameData[184] ;
  wire \FrameData[185] ;
  wire \FrameData[186] ;
  wire \FrameData[187] ;
  wire \FrameData[188] ;
  wire \FrameData[189] ;
  wire \FrameData[190] ;
  wire \FrameData[191] ;
  wire \FrameData[192] ;
  wire \FrameData[193] ;
  wire \FrameData[194] ;
  wire \FrameData[195] ;
  wire \FrameData[196] ;
  wire \FrameData[197] ;
  wire \FrameData[198] ;
  wire \FrameData[199] ;
  wire \FrameData[200] ;
  wire \FrameData[201] ;
  wire \FrameData[202] ;
  wire \FrameData[203] ;
  wire \FrameData[204] ;
  wire \FrameData[205] ;
  wire \FrameData[206] ;
  wire \FrameData[207] ;
  wire \FrameData[208] ;
  wire \FrameData[209] ;
  wire \FrameData[210] ;
  wire \FrameData[211] ;
  wire \FrameData[212] ;
  wire \FrameData[213] ;
  wire \FrameData[214] ;
  wire \FrameData[215] ;
  wire \FrameData[216] ;
  wire \FrameData[217] ;
  wire \FrameData[218] ;
  wire \FrameData[219] ;
  wire \FrameData[220] ;
  wire \FrameData[221] ;
  wire \FrameData[222] ;
  wire \FrameData[223] ;
  wire \FrameData[224] ;
  wire \FrameData[225] ;
  wire \FrameData[226] ;
  wire \FrameData[227] ;
  wire \FrameData[228] ;
  wire \FrameData[229] ;
  wire \FrameData[230] ;
  wire \FrameData[231] ;
  wire \FrameData[232] ;
  wire \FrameData[233] ;
  wire \FrameData[234] ;
  wire \FrameData[235] ;
  wire \FrameData[236] ;
  wire \FrameData[237] ;
  wire \FrameData[238] ;
  wire \FrameData[239] ;
  wire \FrameData[240] ;
  wire \FrameData[241] ;
  wire \FrameData[242] ;
  wire \FrameData[243] ;
  wire \FrameData[244] ;
  wire \FrameData[245] ;
  wire \FrameData[246] ;
  wire \FrameData[247] ;
  wire \FrameData[248] ;
  wire \FrameData[249] ;
  wire \FrameData[250] ;
  wire \FrameData[251] ;
  wire \FrameData[252] ;
  wire \FrameData[253] ;
  wire \FrameData[254] ;
  wire \FrameData[255] ;
  wire \FrameData[256] ;
  wire \FrameData[257] ;
  wire \FrameData[258] ;
  wire \FrameData[259] ;
  wire \FrameData[260] ;
  wire \FrameData[261] ;
  wire \FrameData[262] ;
  wire \FrameData[263] ;
  wire \FrameData[264] ;
  wire \FrameData[265] ;
  wire \FrameData[266] ;
  wire \FrameData[267] ;
  wire \FrameData[268] ;
  wire \FrameData[269] ;
  wire \FrameData[270] ;
  wire \FrameData[271] ;
  wire \FrameData[272] ;
  wire \FrameData[273] ;
  wire \FrameData[274] ;
  wire \FrameData[275] ;
  wire \FrameData[276] ;
  wire \FrameData[277] ;
  wire \FrameData[278] ;
  wire \FrameData[279] ;
  wire \FrameData[280] ;
  wire \FrameData[281] ;
  wire \FrameData[282] ;
  wire \FrameData[283] ;
  wire \FrameData[284] ;
  wire \FrameData[285] ;
  wire \FrameData[286] ;
  wire \FrameData[287] ;
  wire \FrameData[288] ;
  wire \FrameData[289] ;
  wire \FrameData[290] ;
  wire \FrameData[291] ;
  wire \FrameData[292] ;
  wire \FrameData[293] ;
  wire \FrameData[294] ;
  wire \FrameData[295] ;
  wire \FrameData[296] ;
  wire \FrameData[297] ;
  wire \FrameData[298] ;
  wire \FrameData[299] ;
  wire \FrameData[300] ;
  wire \FrameData[301] ;
  wire \FrameData[302] ;
  wire \FrameData[303] ;
  wire \FrameData[304] ;
  wire \FrameData[305] ;
  wire \FrameData[306] ;
  wire \FrameData[307] ;
  wire \FrameData[308] ;
  wire \FrameData[309] ;
  wire \FrameData[310] ;
  wire \FrameData[311] ;
  wire \FrameData[312] ;
  wire \FrameData[313] ;
  wire \FrameData[314] ;
  wire \FrameData[315] ;
  wire \FrameData[316] ;
  wire \FrameData[317] ;
  wire \FrameData[318] ;
  wire \FrameData[319] ;
  wire \FrameData[320] ;
  wire \FrameData[321] ;
  wire \FrameData[322] ;
  wire \FrameData[323] ;
  wire \FrameData[324] ;
  wire \FrameData[325] ;
  wire \FrameData[326] ;
  wire \FrameData[327] ;
  wire \FrameData[328] ;
  wire \FrameData[329] ;
  wire \FrameData[32] ;
  wire \FrameData[330] ;
  wire \FrameData[331] ;
  wire \FrameData[332] ;
  wire \FrameData[333] ;
  wire \FrameData[334] ;
  wire \FrameData[335] ;
  wire \FrameData[336] ;
  wire \FrameData[337] ;
  wire \FrameData[338] ;
  wire \FrameData[339] ;
  wire \FrameData[33] ;
  wire \FrameData[340] ;
  wire \FrameData[341] ;
  wire \FrameData[342] ;
  wire \FrameData[343] ;
  wire \FrameData[344] ;
  wire \FrameData[345] ;
  wire \FrameData[346] ;
  wire \FrameData[347] ;
  wire \FrameData[348] ;
  wire \FrameData[349] ;
  wire \FrameData[34] ;
  wire \FrameData[350] ;
  wire \FrameData[351] ;
  wire \FrameData[352] ;
  wire \FrameData[353] ;
  wire \FrameData[354] ;
  wire \FrameData[355] ;
  wire \FrameData[356] ;
  wire \FrameData[357] ;
  wire \FrameData[358] ;
  wire \FrameData[359] ;
  wire \FrameData[35] ;
  wire \FrameData[360] ;
  wire \FrameData[361] ;
  wire \FrameData[362] ;
  wire \FrameData[363] ;
  wire \FrameData[364] ;
  wire \FrameData[365] ;
  wire \FrameData[366] ;
  wire \FrameData[367] ;
  wire \FrameData[368] ;
  wire \FrameData[369] ;
  wire \FrameData[36] ;
  wire \FrameData[370] ;
  wire \FrameData[371] ;
  wire \FrameData[372] ;
  wire \FrameData[373] ;
  wire \FrameData[374] ;
  wire \FrameData[375] ;
  wire \FrameData[376] ;
  wire \FrameData[377] ;
  wire \FrameData[378] ;
  wire \FrameData[379] ;
  wire \FrameData[37] ;
  wire \FrameData[380] ;
  wire \FrameData[381] ;
  wire \FrameData[382] ;
  wire \FrameData[383] ;
  wire \FrameData[384] ;
  wire \FrameData[385] ;
  wire \FrameData[386] ;
  wire \FrameData[387] ;
  wire \FrameData[388] ;
  wire \FrameData[389] ;
  wire \FrameData[38] ;
  wire \FrameData[390] ;
  wire \FrameData[391] ;
  wire \FrameData[392] ;
  wire \FrameData[393] ;
  wire \FrameData[394] ;
  wire \FrameData[395] ;
  wire \FrameData[396] ;
  wire \FrameData[397] ;
  wire \FrameData[398] ;
  wire \FrameData[399] ;
  wire \FrameData[39] ;
  wire \FrameData[400] ;
  wire \FrameData[401] ;
  wire \FrameData[402] ;
  wire \FrameData[403] ;
  wire \FrameData[404] ;
  wire \FrameData[405] ;
  wire \FrameData[406] ;
  wire \FrameData[407] ;
  wire \FrameData[408] ;
  wire \FrameData[409] ;
  wire \FrameData[40] ;
  wire \FrameData[410] ;
  wire \FrameData[411] ;
  wire \FrameData[412] ;
  wire \FrameData[413] ;
  wire \FrameData[414] ;
  wire \FrameData[415] ;
  wire \FrameData[416] ;
  wire \FrameData[417] ;
  wire \FrameData[418] ;
  wire \FrameData[419] ;
  wire \FrameData[41] ;
  wire \FrameData[420] ;
  wire \FrameData[421] ;
  wire \FrameData[422] ;
  wire \FrameData[423] ;
  wire \FrameData[424] ;
  wire \FrameData[425] ;
  wire \FrameData[426] ;
  wire \FrameData[427] ;
  wire \FrameData[428] ;
  wire \FrameData[429] ;
  wire \FrameData[42] ;
  wire \FrameData[430] ;
  wire \FrameData[431] ;
  wire \FrameData[432] ;
  wire \FrameData[433] ;
  wire \FrameData[434] ;
  wire \FrameData[435] ;
  wire \FrameData[436] ;
  wire \FrameData[437] ;
  wire \FrameData[438] ;
  wire \FrameData[439] ;
  wire \FrameData[43] ;
  wire \FrameData[440] ;
  wire \FrameData[441] ;
  wire \FrameData[442] ;
  wire \FrameData[443] ;
  wire \FrameData[444] ;
  wire \FrameData[445] ;
  wire \FrameData[446] ;
  wire \FrameData[447] ;
  wire \FrameData[448] ;
  wire \FrameData[449] ;
  wire \FrameData[44] ;
  wire \FrameData[450] ;
  wire \FrameData[451] ;
  wire \FrameData[452] ;
  wire \FrameData[453] ;
  wire \FrameData[454] ;
  wire \FrameData[455] ;
  wire \FrameData[456] ;
  wire \FrameData[457] ;
  wire \FrameData[458] ;
  wire \FrameData[459] ;
  wire \FrameData[45] ;
  wire \FrameData[460] ;
  wire \FrameData[461] ;
  wire \FrameData[462] ;
  wire \FrameData[463] ;
  wire \FrameData[464] ;
  wire \FrameData[465] ;
  wire \FrameData[466] ;
  wire \FrameData[467] ;
  wire \FrameData[468] ;
  wire \FrameData[469] ;
  wire \FrameData[46] ;
  wire \FrameData[470] ;
  wire \FrameData[471] ;
  wire \FrameData[472] ;
  wire \FrameData[473] ;
  wire \FrameData[474] ;
  wire \FrameData[475] ;
  wire \FrameData[476] ;
  wire \FrameData[477] ;
  wire \FrameData[478] ;
  wire \FrameData[479] ;
  wire \FrameData[47] ;
  wire \FrameData[48] ;
  wire \FrameData[49] ;
  wire \FrameData[50] ;
  wire \FrameData[51] ;
  wire \FrameData[52] ;
  wire \FrameData[53] ;
  wire \FrameData[54] ;
  wire \FrameData[55] ;
  wire \FrameData[56] ;
  wire \FrameData[57] ;
  wire \FrameData[58] ;
  wire \FrameData[59] ;
  wire \FrameData[60] ;
  wire \FrameData[61] ;
  wire \FrameData[62] ;
  wire \FrameData[63] ;
  wire \FrameData[64] ;
  wire \FrameData[65] ;
  wire \FrameData[66] ;
  wire \FrameData[67] ;
  wire \FrameData[68] ;
  wire \FrameData[69] ;
  wire \FrameData[70] ;
  wire \FrameData[71] ;
  wire \FrameData[72] ;
  wire \FrameData[73] ;
  wire \FrameData[74] ;
  wire \FrameData[75] ;
  wire \FrameData[76] ;
  wire \FrameData[77] ;
  wire \FrameData[78] ;
  wire \FrameData[79] ;
  wire \FrameData[80] ;
  wire \FrameData[81] ;
  wire \FrameData[82] ;
  wire \FrameData[83] ;
  wire \FrameData[84] ;
  wire \FrameData[85] ;
  wire \FrameData[86] ;
  wire \FrameData[87] ;
  wire \FrameData[88] ;
  wire \FrameData[89] ;
  wire \FrameData[90] ;
  wire \FrameData[91] ;
  wire \FrameData[92] ;
  wire \FrameData[93] ;
  wire \FrameData[94] ;
  wire \FrameData[95] ;
  wire \FrameData[96] ;
  wire \FrameData[97] ;
  wire \FrameData[98] ;
  wire \FrameData[99] ;
  wire \FrameSelect[0] ;
  wire \FrameSelect[100] ;
  wire \FrameSelect[101] ;
  wire \FrameSelect[102] ;
  wire \FrameSelect[103] ;
  wire \FrameSelect[104] ;
  wire \FrameSelect[105] ;
  wire \FrameSelect[106] ;
  wire \FrameSelect[107] ;
  wire \FrameSelect[108] ;
  wire \FrameSelect[109] ;
  wire \FrameSelect[10] ;
  wire \FrameSelect[110] ;
  wire \FrameSelect[111] ;
  wire \FrameSelect[112] ;
  wire \FrameSelect[113] ;
  wire \FrameSelect[114] ;
  wire \FrameSelect[115] ;
  wire \FrameSelect[116] ;
  wire \FrameSelect[117] ;
  wire \FrameSelect[118] ;
  wire \FrameSelect[119] ;
  wire \FrameSelect[11] ;
  wire \FrameSelect[120] ;
  wire \FrameSelect[121] ;
  wire \FrameSelect[122] ;
  wire \FrameSelect[123] ;
  wire \FrameSelect[124] ;
  wire \FrameSelect[125] ;
  wire \FrameSelect[126] ;
  wire \FrameSelect[127] ;
  wire \FrameSelect[128] ;
  wire \FrameSelect[129] ;
  wire \FrameSelect[12] ;
  wire \FrameSelect[130] ;
  wire \FrameSelect[131] ;
  wire \FrameSelect[132] ;
  wire \FrameSelect[133] ;
  wire \FrameSelect[134] ;
  wire \FrameSelect[135] ;
  wire \FrameSelect[136] ;
  wire \FrameSelect[137] ;
  wire \FrameSelect[138] ;
  wire \FrameSelect[139] ;
  wire \FrameSelect[13] ;
  wire \FrameSelect[140] ;
  wire \FrameSelect[141] ;
  wire \FrameSelect[142] ;
  wire \FrameSelect[143] ;
  wire \FrameSelect[144] ;
  wire \FrameSelect[145] ;
  wire \FrameSelect[146] ;
  wire \FrameSelect[147] ;
  wire \FrameSelect[148] ;
  wire \FrameSelect[149] ;
  wire \FrameSelect[14] ;
  wire \FrameSelect[150] ;
  wire \FrameSelect[151] ;
  wire \FrameSelect[152] ;
  wire \FrameSelect[153] ;
  wire \FrameSelect[154] ;
  wire \FrameSelect[155] ;
  wire \FrameSelect[156] ;
  wire \FrameSelect[157] ;
  wire \FrameSelect[158] ;
  wire \FrameSelect[159] ;
  wire \FrameSelect[15] ;
  wire \FrameSelect[160] ;
  wire \FrameSelect[161] ;
  wire \FrameSelect[162] ;
  wire \FrameSelect[163] ;
  wire \FrameSelect[164] ;
  wire \FrameSelect[165] ;
  wire \FrameSelect[166] ;
  wire \FrameSelect[167] ;
  wire \FrameSelect[168] ;
  wire \FrameSelect[169] ;
  wire \FrameSelect[16] ;
  wire \FrameSelect[170] ;
  wire \FrameSelect[171] ;
  wire \FrameSelect[172] ;
  wire \FrameSelect[173] ;
  wire \FrameSelect[174] ;
  wire \FrameSelect[175] ;
  wire \FrameSelect[176] ;
  wire \FrameSelect[177] ;
  wire \FrameSelect[178] ;
  wire \FrameSelect[179] ;
  wire \FrameSelect[17] ;
  wire \FrameSelect[180] ;
  wire \FrameSelect[181] ;
  wire \FrameSelect[182] ;
  wire \FrameSelect[183] ;
  wire \FrameSelect[184] ;
  wire \FrameSelect[185] ;
  wire \FrameSelect[186] ;
  wire \FrameSelect[187] ;
  wire \FrameSelect[188] ;
  wire \FrameSelect[189] ;
  wire \FrameSelect[18] ;
  wire \FrameSelect[190] ;
  wire \FrameSelect[191] ;
  wire \FrameSelect[192] ;
  wire \FrameSelect[193] ;
  wire \FrameSelect[194] ;
  wire \FrameSelect[195] ;
  wire \FrameSelect[196] ;
  wire \FrameSelect[197] ;
  wire \FrameSelect[198] ;
  wire \FrameSelect[199] ;
  wire \FrameSelect[19] ;
  wire \FrameSelect[1] ;
  wire \FrameSelect[200] ;
  wire \FrameSelect[201] ;
  wire \FrameSelect[202] ;
  wire \FrameSelect[203] ;
  wire \FrameSelect[204] ;
  wire \FrameSelect[205] ;
  wire \FrameSelect[206] ;
  wire \FrameSelect[207] ;
  wire \FrameSelect[208] ;
  wire \FrameSelect[209] ;
  wire \FrameSelect[20] ;
  wire \FrameSelect[210] ;
  wire \FrameSelect[211] ;
  wire \FrameSelect[212] ;
  wire \FrameSelect[213] ;
  wire \FrameSelect[214] ;
  wire \FrameSelect[215] ;
  wire \FrameSelect[216] ;
  wire \FrameSelect[217] ;
  wire \FrameSelect[218] ;
  wire \FrameSelect[219] ;
  wire \FrameSelect[21] ;
  wire \FrameSelect[220] ;
  wire \FrameSelect[221] ;
  wire \FrameSelect[222] ;
  wire \FrameSelect[223] ;
  wire \FrameSelect[224] ;
  wire \FrameSelect[225] ;
  wire \FrameSelect[226] ;
  wire \FrameSelect[227] ;
  wire \FrameSelect[228] ;
  wire \FrameSelect[229] ;
  wire \FrameSelect[22] ;
  wire \FrameSelect[230] ;
  wire \FrameSelect[231] ;
  wire \FrameSelect[232] ;
  wire \FrameSelect[233] ;
  wire \FrameSelect[234] ;
  wire \FrameSelect[235] ;
  wire \FrameSelect[236] ;
  wire \FrameSelect[237] ;
  wire \FrameSelect[238] ;
  wire \FrameSelect[239] ;
  wire \FrameSelect[23] ;
  wire \FrameSelect[240] ;
  wire \FrameSelect[241] ;
  wire \FrameSelect[242] ;
  wire \FrameSelect[243] ;
  wire \FrameSelect[244] ;
  wire \FrameSelect[245] ;
  wire \FrameSelect[246] ;
  wire \FrameSelect[247] ;
  wire \FrameSelect[248] ;
  wire \FrameSelect[249] ;
  wire \FrameSelect[24] ;
  wire \FrameSelect[250] ;
  wire \FrameSelect[251] ;
  wire \FrameSelect[252] ;
  wire \FrameSelect[253] ;
  wire \FrameSelect[254] ;
  wire \FrameSelect[255] ;
  wire \FrameSelect[256] ;
  wire \FrameSelect[257] ;
  wire \FrameSelect[258] ;
  wire \FrameSelect[259] ;
  wire \FrameSelect[25] ;
  wire \FrameSelect[260] ;
  wire \FrameSelect[261] ;
  wire \FrameSelect[262] ;
  wire \FrameSelect[263] ;
  wire \FrameSelect[264] ;
  wire \FrameSelect[265] ;
  wire \FrameSelect[266] ;
  wire \FrameSelect[267] ;
  wire \FrameSelect[268] ;
  wire \FrameSelect[269] ;
  wire \FrameSelect[26] ;
  wire \FrameSelect[270] ;
  wire \FrameSelect[271] ;
  wire \FrameSelect[272] ;
  wire \FrameSelect[273] ;
  wire \FrameSelect[274] ;
  wire \FrameSelect[275] ;
  wire \FrameSelect[276] ;
  wire \FrameSelect[277] ;
  wire \FrameSelect[278] ;
  wire \FrameSelect[279] ;
  wire \FrameSelect[27] ;
  wire \FrameSelect[280] ;
  wire \FrameSelect[281] ;
  wire \FrameSelect[282] ;
  wire \FrameSelect[283] ;
  wire \FrameSelect[284] ;
  wire \FrameSelect[285] ;
  wire \FrameSelect[286] ;
  wire \FrameSelect[287] ;
  wire \FrameSelect[288] ;
  wire \FrameSelect[289] ;
  wire \FrameSelect[28] ;
  wire \FrameSelect[290] ;
  wire \FrameSelect[291] ;
  wire \FrameSelect[292] ;
  wire \FrameSelect[293] ;
  wire \FrameSelect[294] ;
  wire \FrameSelect[295] ;
  wire \FrameSelect[296] ;
  wire \FrameSelect[297] ;
  wire \FrameSelect[298] ;
  wire \FrameSelect[299] ;
  wire \FrameSelect[29] ;
  wire \FrameSelect[2] ;
  wire \FrameSelect[30] ;
  wire \FrameSelect[31] ;
  wire \FrameSelect[32] ;
  wire \FrameSelect[33] ;
  wire \FrameSelect[34] ;
  wire \FrameSelect[35] ;
  wire \FrameSelect[36] ;
  wire \FrameSelect[37] ;
  wire \FrameSelect[38] ;
  wire \FrameSelect[39] ;
  wire \FrameSelect[3] ;
  wire \FrameSelect[40] ;
  wire \FrameSelect[41] ;
  wire \FrameSelect[42] ;
  wire \FrameSelect[43] ;
  wire \FrameSelect[44] ;
  wire \FrameSelect[45] ;
  wire \FrameSelect[46] ;
  wire \FrameSelect[47] ;
  wire \FrameSelect[48] ;
  wire \FrameSelect[49] ;
  wire \FrameSelect[4] ;
  wire \FrameSelect[50] ;
  wire \FrameSelect[51] ;
  wire \FrameSelect[52] ;
  wire \FrameSelect[53] ;
  wire \FrameSelect[54] ;
  wire \FrameSelect[55] ;
  wire \FrameSelect[56] ;
  wire \FrameSelect[57] ;
  wire \FrameSelect[58] ;
  wire \FrameSelect[59] ;
  wire \FrameSelect[5] ;
  wire \FrameSelect[60] ;
  wire \FrameSelect[61] ;
  wire \FrameSelect[62] ;
  wire \FrameSelect[63] ;
  wire \FrameSelect[64] ;
  wire \FrameSelect[65] ;
  wire \FrameSelect[66] ;
  wire \FrameSelect[67] ;
  wire \FrameSelect[68] ;
  wire \FrameSelect[69] ;
  wire \FrameSelect[6] ;
  wire \FrameSelect[70] ;
  wire \FrameSelect[71] ;
  wire \FrameSelect[72] ;
  wire \FrameSelect[73] ;
  wire \FrameSelect[74] ;
  wire \FrameSelect[75] ;
  wire \FrameSelect[76] ;
  wire \FrameSelect[77] ;
  wire \FrameSelect[78] ;
  wire \FrameSelect[79] ;
  wire \FrameSelect[7] ;
  wire \FrameSelect[80] ;
  wire \FrameSelect[81] ;
  wire \FrameSelect[82] ;
  wire \FrameSelect[83] ;
  wire \FrameSelect[84] ;
  wire \FrameSelect[85] ;
  wire \FrameSelect[86] ;
  wire \FrameSelect[87] ;
  wire \FrameSelect[88] ;
  wire \FrameSelect[89] ;
  wire \FrameSelect[8] ;
  wire \FrameSelect[90] ;
  wire \FrameSelect[91] ;
  wire \FrameSelect[92] ;
  wire \FrameSelect[93] ;
  wire \FrameSelect[94] ;
  wire \FrameSelect[95] ;
  wire \FrameSelect[96] ;
  wire \FrameSelect[97] ;
  wire \FrameSelect[98] ;
  wire \FrameSelect[99] ;
  wire \FrameSelect[9] ;
  wire \LocalWriteData[0] ;
  wire \LocalWriteData[10] ;
  wire \LocalWriteData[11] ;
  wire \LocalWriteData[12] ;
  wire \LocalWriteData[13] ;
  wire \LocalWriteData[14] ;
  wire \LocalWriteData[15] ;
  wire \LocalWriteData[16] ;
  wire \LocalWriteData[17] ;
  wire \LocalWriteData[18] ;
  wire \LocalWriteData[19] ;
  wire \LocalWriteData[1] ;
  wire \LocalWriteData[20] ;
  wire \LocalWriteData[21] ;
  wire \LocalWriteData[22] ;
  wire \LocalWriteData[23] ;
  wire \LocalWriteData[24] ;
  wire \LocalWriteData[25] ;
  wire \LocalWriteData[26] ;
  wire \LocalWriteData[27] ;
  wire \LocalWriteData[28] ;
  wire \LocalWriteData[29] ;
  wire \LocalWriteData[2] ;
  wire \LocalWriteData[30] ;
  wire \LocalWriteData[31] ;
  wire \LocalWriteData[3] ;
  wire \LocalWriteData[4] ;
  wire \LocalWriteData[5] ;
  wire \LocalWriteData[6] ;
  wire \LocalWriteData[7] ;
  wire \LocalWriteData[8] ;
  wire \LocalWriteData[9] ;
  wire LocalWriteStrobe;
  wire LongFrameStrobe;
  wire ReceiveLED;
  wire \RowSelect[0] ;
  wire \RowSelect[1] ;
  wire \RowSelect[2] ;
  wire \RowSelect[3] ;
  wire \RowSelect[4] ;
  wire \SelfWriteData[0] ;
  wire \SelfWriteData[10] ;
  wire \SelfWriteData[11] ;
  wire \SelfWriteData[12] ;
  wire \SelfWriteData[13] ;
  wire \SelfWriteData[14] ;
  wire \SelfWriteData[15] ;
  wire \SelfWriteData[16] ;
  wire \SelfWriteData[17] ;
  wire \SelfWriteData[18] ;
  wire \SelfWriteData[19] ;
  wire \SelfWriteData[1] ;
  wire \SelfWriteData[20] ;
  wire \SelfWriteData[21] ;
  wire \SelfWriteData[22] ;
  wire \SelfWriteData[23] ;
  wire \SelfWriteData[24] ;
  wire \SelfWriteData[25] ;
  wire \SelfWriteData[26] ;
  wire \SelfWriteData[27] ;
  wire \SelfWriteData[28] ;
  wire \SelfWriteData[29] ;
  wire \SelfWriteData[2] ;
  wire \SelfWriteData[30] ;
  wire \SelfWriteData[31] ;
  wire \SelfWriteData[3] ;
  wire \SelfWriteData[4] ;
  wire \SelfWriteData[5] ;
  wire \SelfWriteData[6] ;
  wire \SelfWriteData[7] ;
  wire \SelfWriteData[8] ;
  wire \SelfWriteData[9] ;
  wire SelfWriteStrobe;
  wire \W_OPA[0] ;
  wire \W_OPA[1] ;
  wire \W_OPA[2] ;
  wire \W_OPA[35] ;
  wire \W_OPB[0] ;
  wire \W_OPB[10] ;
  wire \W_OPB[11] ;
  wire \W_OPB[12] ;
  wire \W_OPB[13] ;
  wire \W_OPB[14] ;
  wire \W_OPB[15] ;
  wire \W_OPB[16] ;
  wire \W_OPB[17] ;
  wire \W_OPB[18] ;
  wire \W_OPB[19] ;
  wire \W_OPB[1] ;
  wire \W_OPB[20] ;
  wire \W_OPB[21] ;
  wire \W_OPB[22] ;
  wire \W_OPB[23] ;
  wire \W_OPB[24] ;
  wire \W_OPB[25] ;
  wire \W_OPB[26] ;
  wire \W_OPB[27] ;
  wire \W_OPB[28] ;
  wire \W_OPB[29] ;
  wire \W_OPB[2] ;
  wire \W_OPB[30] ;
  wire \W_OPB[31] ;
  wire \W_OPB[32] ;
  wire \W_OPB[33] ;
  wire \W_OPB[34] ;
  wire \W_OPB[35] ;
  wire \W_OPB[3] ;
  wire \W_OPB[4] ;
  wire \W_OPB[5] ;
  wire \W_OPB[6] ;
  wire \W_OPB[7] ;
  wire \W_OPB[8] ;
  wire \W_OPB[9] ;
  wire \W_RES0[0] ;
  wire \W_RES0[10] ;
  wire \W_RES0[11] ;
  wire \W_RES0[12] ;
  wire \W_RES0[13] ;
  wire \W_RES0[14] ;
  wire \W_RES0[15] ;
  wire \W_RES0[16] ;
  wire \W_RES0[17] ;
  wire \W_RES0[18] ;
  wire \W_RES0[19] ;
  wire \W_RES0[1] ;
  wire \W_RES0[20] ;
  wire \W_RES0[21] ;
  wire \W_RES0[22] ;
  wire \W_RES0[23] ;
  wire \W_RES0[24] ;
  wire \W_RES0[25] ;
  wire \W_RES0[26] ;
  wire \W_RES0[27] ;
  wire \W_RES0[28] ;
  wire \W_RES0[29] ;
  wire \W_RES0[2] ;
  wire \W_RES0[30] ;
  wire \W_RES0[31] ;
  wire \W_RES0[32] ;
  wire \W_RES0[33] ;
  wire \W_RES0[34] ;
  wire \W_RES0[35] ;
  wire \W_RES0[3] ;
  wire \W_RES0[4] ;
  wire \W_RES0[5] ;
  wire \W_RES0[6] ;
  wire \W_RES0[7] ;
  wire \W_RES0[8] ;
  wire \W_RES0[9] ;
  wire \W_RES1[0] ;
  wire \W_RES1[10] ;
  wire \W_RES1[11] ;
  wire \W_RES1[12] ;
  wire \W_RES1[13] ;
  wire \W_RES1[14] ;
  wire \W_RES1[15] ;
  wire \W_RES1[16] ;
  wire \W_RES1[17] ;
  wire \W_RES1[18] ;
  wire \W_RES1[19] ;
  wire \W_RES1[1] ;
  wire \W_RES1[20] ;
  wire \W_RES1[21] ;
  wire \W_RES1[22] ;
  wire \W_RES1[23] ;
  wire \W_RES1[24] ;
  wire \W_RES1[25] ;
  wire \W_RES1[26] ;
  wire \W_RES1[27] ;
  wire \W_RES1[28] ;
  wire \W_RES1[29] ;
  wire \W_RES1[2] ;
  wire \W_RES1[30] ;
  wire \W_RES1[31] ;
  wire \W_RES1[32] ;
  wire \W_RES1[33] ;
  wire \W_RES1[34] ;
  wire \W_RES1[35] ;
  wire \W_RES1[3] ;
  wire \W_RES1[4] ;
  wire \W_RES1[5] ;
  wire \W_RES1[6] ;
  wire \W_RES1[7] ;
  wire \W_RES1[8] ;
  wire \W_RES1[9] ;
  wire \W_RES2[0] ;
  wire \W_RES2[10] ;
  wire \W_RES2[11] ;
  wire \W_RES2[12] ;
  wire \W_RES2[13] ;
  wire \W_RES2[14] ;
  wire \W_RES2[15] ;
  wire \W_RES2[16] ;
  wire \W_RES2[17] ;
  wire \W_RES2[18] ;
  wire \W_RES2[19] ;
  wire \W_RES2[1] ;
  wire \W_RES2[20] ;
  wire \W_RES2[21] ;
  wire \W_RES2[22] ;
  wire \W_RES2[23] ;
  wire \W_RES2[24] ;
  wire \W_RES2[25] ;
  wire \W_RES2[26] ;
  wire \W_RES2[27] ;
  wire \W_RES2[28] ;
  wire \W_RES2[29] ;
  wire \W_RES2[2] ;
  wire \W_RES2[30] ;
  wire \W_RES2[31] ;
  wire \W_RES2[32] ;
  wire \W_RES2[33] ;
  wire \W_RES2[34] ;
  wire \W_RES2[35] ;
  wire \W_RES2[3] ;
  wire \W_RES2[4] ;
  wire \W_RES2[5] ;
  wire \W_RES2[6] ;
  wire \W_RES2[7] ;
  wire \W_RES2[8] ;
  wire \W_RES2[9] ;
  wire debug_req_1;
  wire debug_req_2;
  wire fetch_enable_1;
  wire fetch_enable_2;
  input [37:0] io_in;
  output [37:0] io_oeb;
  output [37:0] io_out;
  input [3:0] la_data_in;
  output [2:0] la_data_out;
  input user_clock2;
  input wb_clk_i;
  input wb_rst_i;
  output wbs_ack_o;
  input [31:0] wbs_adr_i;
  input wbs_cyc_i;
  input [31:0] wbs_dat_i;
  output [31:0] wbs_dat_o;
  input [3:0] wbs_sel_i;
  input wbs_stb_i;
  input wbs_we_i;
  sky130_fd_sc_hd__conb_1 _155_ (
    .HI(_011_)
  );
  sky130_fd_sc_hd__conb_1 _156_ (
    .HI(_012_)
  );
  sky130_fd_sc_hd__conb_1 _157_ (
    .HI(_013_)
  );
  sky130_fd_sc_hd__conb_1 _158_ (
    .HI(_014_)
  );
  sky130_fd_sc_hd__conb_1 _159_ (
    .HI(_015_)
  );
  sky130_fd_sc_hd__conb_1 _160_ (
    .HI(_016_)
  );
  sky130_fd_sc_hd__conb_1 _161_ (
    .HI(_017_)
  );
  sky130_fd_sc_hd__conb_1 _162_ (
    .HI(_018_)
  );
  sky130_fd_sc_hd__conb_1 _163_ (
    .HI(_019_)
  );
  sky130_fd_sc_hd__conb_1 _164_ (
    .HI(_020_)
  );
  sky130_fd_sc_hd__conb_1 _165_ (
    .HI(_021_)
  );
  sky130_fd_sc_hd__conb_1 _166_ (
    .HI(_022_)
  );
  sky130_fd_sc_hd__conb_1 _167_ (
    .HI(_023_)
  );
  sky130_fd_sc_hd__conb_1 _168_ (
    .HI(_024_)
  );
  sky130_fd_sc_hd__conb_1 _169_ (
    .HI(_025_)
  );
  sky130_fd_sc_hd__conb_1 _170_ (
    .HI(_026_)
  );
  sky130_fd_sc_hd__conb_1 _171_ (
    .HI(_027_)
  );
  sky130_fd_sc_hd__conb_1 _172_ (
    .HI(_028_)
  );
  sky130_fd_sc_hd__conb_1 _173_ (
    .HI(_029_)
  );
  sky130_fd_sc_hd__conb_1 _174_ (
    .HI(_030_)
  );
  sky130_fd_sc_hd__conb_1 _175_ (
    .HI(_031_)
  );
  sky130_fd_sc_hd__conb_1 _176_ (
    .HI(_032_)
  );
  sky130_fd_sc_hd__conb_1 _177_ (
    .HI(_033_)
  );
  sky130_fd_sc_hd__conb_1 _178_ (
    .HI(_034_)
  );
  sky130_fd_sc_hd__conb_1 _179_ (
    .HI(_035_)
  );
  sky130_fd_sc_hd__conb_1 _180_ (
    .HI(_036_)
  );
  sky130_fd_sc_hd__conb_1 _181_ (
    .HI(io_oeb[0])
  );
  sky130_fd_sc_hd__conb_1 _182_ (
    .HI(io_oeb[1])
  );
  sky130_fd_sc_hd__conb_1 _183_ (
    .HI(io_oeb[2])
  );
  sky130_fd_sc_hd__conb_1 _184_ (
    .HI(io_oeb[3])
  );
  sky130_fd_sc_hd__conb_1 _185_ (
    .HI(io_oeb[4])
  );
  sky130_fd_sc_hd__conb_1 _186_ (
    .HI(io_oeb[5])
  );
  sky130_fd_sc_hd__conb_1 _187_ (
    .HI(io_oeb[7])
  );
  sky130_fd_sc_hd__conb_1 _188_ (
    .HI(io_oeb[8])
  );
  sky130_fd_sc_hd__conb_1 _189_ (
    .HI(io_oeb[9])
  );
  sky130_fd_sc_hd__conb_1 _190_ (
    .HI(io_oeb[10])
  );
  sky130_fd_sc_hd__conb_1 _191_ (
    .HI(io_oeb[11])
  );
  sky130_fd_sc_hd__conb_1 _192_ (
    .HI(io_oeb[12])
  );
  sky130_fd_sc_hd__conb_1 _193_ (
    .HI(io_oeb[14])
  );
  sky130_fd_sc_hd__conb_1 _194_ (
    .LO(_037_)
  );
  sky130_fd_sc_hd__conb_1 _195_ (
    .LO(_038_)
  );
  sky130_fd_sc_hd__conb_1 _196_ (
    .LO(_039_)
  );
  sky130_fd_sc_hd__conb_1 _197_ (
    .LO(_040_)
  );
  sky130_fd_sc_hd__conb_1 _198_ (
    .LO(_041_)
  );
  sky130_fd_sc_hd__conb_1 _199_ (
    .LO(_042_)
  );
  sky130_fd_sc_hd__conb_1 _200_ (
    .LO(_043_)
  );
  sky130_fd_sc_hd__conb_1 _201_ (
    .LO(_044_)
  );
  sky130_fd_sc_hd__conb_1 _202_ (
    .LO(_045_)
  );
  sky130_fd_sc_hd__conb_1 _203_ (
    .LO(_046_)
  );
  sky130_fd_sc_hd__conb_1 _204_ (
    .LO(_047_)
  );
  sky130_fd_sc_hd__conb_1 _205_ (
    .LO(_048_)
  );
  sky130_fd_sc_hd__conb_1 _206_ (
    .LO(_049_)
  );
  sky130_fd_sc_hd__conb_1 _207_ (
    .LO(_050_)
  );
  sky130_fd_sc_hd__conb_1 _208_ (
    .LO(_051_)
  );
  sky130_fd_sc_hd__conb_1 _209_ (
    .LO(_052_)
  );
  sky130_fd_sc_hd__conb_1 _210_ (
    .LO(_053_)
  );
  sky130_fd_sc_hd__conb_1 _211_ (
    .LO(_054_)
  );
  sky130_fd_sc_hd__conb_1 _212_ (
    .LO(_055_)
  );
  sky130_fd_sc_hd__conb_1 _213_ (
    .LO(_056_)
  );
  sky130_fd_sc_hd__conb_1 _214_ (
    .LO(_057_)
  );
  sky130_fd_sc_hd__conb_1 _215_ (
    .LO(_058_)
  );
  sky130_fd_sc_hd__conb_1 _216_ (
    .LO(_059_)
  );
  sky130_fd_sc_hd__conb_1 _217_ (
    .LO(_060_)
  );
  sky130_fd_sc_hd__conb_1 _218_ (
    .LO(_061_)
  );
  sky130_fd_sc_hd__conb_1 _219_ (
    .LO(_062_)
  );
  sky130_fd_sc_hd__conb_1 _220_ (
    .LO(_063_)
  );
  sky130_fd_sc_hd__conb_1 _221_ (
    .LO(_064_)
  );
  sky130_fd_sc_hd__conb_1 _222_ (
    .LO(_065_)
  );
  sky130_fd_sc_hd__conb_1 _223_ (
    .LO(_066_)
  );
  sky130_fd_sc_hd__conb_1 _224_ (
    .LO(_067_)
  );
  sky130_fd_sc_hd__conb_1 _225_ (
    .LO(_068_)
  );
  sky130_fd_sc_hd__conb_1 _226_ (
    .LO(_069_)
  );
  sky130_fd_sc_hd__conb_1 _227_ (
    .LO(_070_)
  );
  sky130_fd_sc_hd__conb_1 _228_ (
    .LO(_071_)
  );
  sky130_fd_sc_hd__conb_1 _229_ (
    .LO(_072_)
  );
  sky130_fd_sc_hd__conb_1 _230_ (
    .LO(_073_)
  );
  sky130_fd_sc_hd__conb_1 _231_ (
    .LO(_074_)
  );
  sky130_fd_sc_hd__conb_1 _232_ (
    .LO(_075_)
  );
  sky130_fd_sc_hd__conb_1 _233_ (
    .LO(_076_)
  );
  sky130_fd_sc_hd__conb_1 _234_ (
    .LO(_077_)
  );
  sky130_fd_sc_hd__conb_1 _235_ (
    .LO(_078_)
  );
  sky130_fd_sc_hd__conb_1 _236_ (
    .LO(_079_)
  );
  sky130_fd_sc_hd__conb_1 _237_ (
    .LO(_080_)
  );
  sky130_fd_sc_hd__conb_1 _238_ (
    .LO(_081_)
  );
  sky130_fd_sc_hd__conb_1 _239_ (
    .LO(_082_)
  );
  sky130_fd_sc_hd__conb_1 _240_ (
    .LO(_083_)
  );
  sky130_fd_sc_hd__conb_1 _241_ (
    .LO(_084_)
  );
  sky130_fd_sc_hd__conb_1 _242_ (
    .LO(_085_)
  );
  sky130_fd_sc_hd__conb_1 _243_ (
    .LO(_086_)
  );
  sky130_fd_sc_hd__conb_1 _244_ (
    .LO(_087_)
  );
  sky130_fd_sc_hd__conb_1 _245_ (
    .LO(_088_)
  );
  sky130_fd_sc_hd__conb_1 _246_ (
    .LO(_089_)
  );
  sky130_fd_sc_hd__conb_1 _247_ (
    .LO(_090_)
  );
  sky130_fd_sc_hd__conb_1 _248_ (
    .LO(_091_)
  );
  sky130_fd_sc_hd__conb_1 _249_ (
    .LO(_092_)
  );
  sky130_fd_sc_hd__conb_1 _250_ (
    .LO(_093_)
  );
  sky130_fd_sc_hd__conb_1 _251_ (
    .LO(_094_)
  );
  sky130_fd_sc_hd__conb_1 _252_ (
    .LO(_095_)
  );
  sky130_fd_sc_hd__conb_1 _253_ (
    .LO(_096_)
  );
  sky130_fd_sc_hd__conb_1 _254_ (
    .LO(_097_)
  );
  sky130_fd_sc_hd__conb_1 _255_ (
    .LO(_098_)
  );
  sky130_fd_sc_hd__conb_1 _256_ (
    .LO(_099_)
  );
  sky130_fd_sc_hd__conb_1 _257_ (
    .LO(_100_)
  );
  sky130_fd_sc_hd__conb_1 _258_ (
    .LO(_101_)
  );
  sky130_fd_sc_hd__conb_1 _259_ (
    .LO(_102_)
  );
  sky130_fd_sc_hd__conb_1 _260_ (
    .LO(_103_)
  );
  sky130_fd_sc_hd__conb_1 _261_ (
    .LO(_104_)
  );
  sky130_fd_sc_hd__conb_1 _262_ (
    .LO(_105_)
  );
  sky130_fd_sc_hd__conb_1 _263_ (
    .LO(_106_)
  );
  sky130_fd_sc_hd__conb_1 _264_ (
    .LO(_107_)
  );
  sky130_fd_sc_hd__conb_1 _265_ (
    .LO(_108_)
  );
  sky130_fd_sc_hd__conb_1 _266_ (
    .LO(_109_)
  );
  sky130_fd_sc_hd__conb_1 _267_ (
    .LO(_110_)
  );
  sky130_fd_sc_hd__conb_1 _268_ (
    .LO(_111_)
  );
  sky130_fd_sc_hd__conb_1 _269_ (
    .LO(_112_)
  );
  sky130_fd_sc_hd__conb_1 _270_ (
    .LO(_113_)
  );
  sky130_fd_sc_hd__conb_1 _271_ (
    .LO(_114_)
  );
  sky130_fd_sc_hd__conb_1 _272_ (
    .LO(_115_)
  );
  sky130_fd_sc_hd__conb_1 _273_ (
    .LO(_116_)
  );
  sky130_fd_sc_hd__conb_1 _274_ (
    .LO(_117_)
  );
  sky130_fd_sc_hd__conb_1 _275_ (
    .LO(_118_)
  );
  sky130_fd_sc_hd__conb_1 _276_ (
    .LO(_119_)
  );
  sky130_fd_sc_hd__conb_1 _277_ (
    .LO(_120_)
  );
  sky130_fd_sc_hd__conb_1 _278_ (
    .LO(_121_)
  );
  sky130_fd_sc_hd__conb_1 _279_ (
    .LO(_122_)
  );
  sky130_fd_sc_hd__conb_1 _280_ (
    .LO(_123_)
  );
  sky130_fd_sc_hd__conb_1 _281_ (
    .LO(_124_)
  );
  sky130_fd_sc_hd__conb_1 _282_ (
    .LO(_125_)
  );
  sky130_fd_sc_hd__conb_1 _283_ (
    .LO(_126_)
  );
  sky130_fd_sc_hd__conb_1 _284_ (
    .LO(_127_)
  );
  sky130_fd_sc_hd__conb_1 _285_ (
    .LO(_128_)
  );
  sky130_fd_sc_hd__conb_1 _286_ (
    .LO(_129_)
  );
  sky130_fd_sc_hd__conb_1 _287_ (
    .LO(_130_)
  );
  sky130_fd_sc_hd__conb_1 _288_ (
    .LO(_131_)
  );
  sky130_fd_sc_hd__conb_1 _289_ (
    .LO(_132_)
  );
  sky130_fd_sc_hd__conb_1 _290_ (
    .LO(_133_)
  );
  sky130_fd_sc_hd__conb_1 _291_ (
    .LO(_134_)
  );
  sky130_fd_sc_hd__conb_1 _292_ (
    .LO(_135_)
  );
  sky130_fd_sc_hd__conb_1 _293_ (
    .LO(_136_)
  );
  sky130_fd_sc_hd__conb_1 _294_ (
    .LO(_137_)
  );
  sky130_fd_sc_hd__conb_1 _295_ (
    .LO(_138_)
  );
  sky130_fd_sc_hd__conb_1 _296_ (
    .LO(_139_)
  );
  sky130_fd_sc_hd__conb_1 _297_ (
    .LO(_140_)
  );
  sky130_fd_sc_hd__conb_1 _298_ (
    .LO(_141_)
  );
  sky130_fd_sc_hd__conb_1 _299_ (
    .LO(_142_)
  );
  sky130_fd_sc_hd__conb_1 _300_ (
    .LO(_143_)
  );
  sky130_fd_sc_hd__conb_1 _301_ (
    .LO(_144_)
  );
  sky130_fd_sc_hd__conb_1 _302_ (
    .LO(_145_)
  );
  sky130_fd_sc_hd__conb_1 _303_ (
    .LO(_146_)
  );
  sky130_fd_sc_hd__conb_1 _304_ (
    .LO(_147_)
  );
  sky130_fd_sc_hd__conb_1 _305_ (
    .LO(_148_)
  );
  sky130_fd_sc_hd__conb_1 _306_ (
    .LO(_149_)
  );
  sky130_fd_sc_hd__conb_1 _307_ (
    .LO(_150_)
  );
  sky130_fd_sc_hd__conb_1 _308_ (
    .LO(_151_)
  );
  sky130_fd_sc_hd__conb_1 _309_ (
    .LO(_152_)
  );
  sky130_fd_sc_hd__conb_1 _310_ (
    .LO(_153_)
  );
  sky130_fd_sc_hd__conb_1 _311_ (
    .LO(_154_)
  );
  sky130_fd_sc_hd__conb_1 _312_ (
    .LO(io_oeb[6])
  );
  sky130_fd_sc_hd__conb_1 _313_ (
    .LO(io_oeb[13])
  );
  sky130_fd_sc_hd__conb_1 _314_ (
    .LO(io_oeb[15])
  );
  sky130_fd_sc_hd__conb_1 _315_ (
    .LO(io_oeb[16])
  );
  sky130_fd_sc_hd__conb_1 _316_ (
    .LO(io_oeb[27])
  );
  sky130_fd_sc_hd__conb_1 _317_ (
    .LO(io_oeb[28])
  );
  sky130_fd_sc_hd__conb_1 _318_ (
    .LO(io_oeb[29])
  );
  sky130_fd_sc_hd__conb_1 _319_ (
    .LO(io_oeb[30])
  );
  sky130_fd_sc_hd__conb_1 _320_ (
    .LO(io_oeb[31])
  );
  sky130_fd_sc_hd__conb_1 _321_ (
    .LO(io_oeb[32])
  );
  sky130_fd_sc_hd__conb_1 _322_ (
    .LO(io_oeb[33])
  );
  sky130_fd_sc_hd__conb_1 _323_ (
    .LO(io_oeb[34])
  );
  sky130_fd_sc_hd__conb_1 _324_ (
    .LO(io_oeb[35])
  );
  sky130_fd_sc_hd__conb_1 _325_ (
    .LO(io_oeb[36])
  );
  sky130_fd_sc_hd__conb_1 _326_ (
    .LO(io_oeb[37])
  );
  sky130_fd_sc_hd__conb_1 _327_ (
    .LO(io_out[0])
  );
  sky130_fd_sc_hd__conb_1 _328_ (
    .LO(io_out[1])
  );
  sky130_fd_sc_hd__conb_1 _329_ (
    .LO(io_out[2])
  );
  sky130_fd_sc_hd__conb_1 _330_ (
    .LO(io_out[3])
  );
  sky130_fd_sc_hd__conb_1 _331_ (
    .LO(io_out[4])
  );
  sky130_fd_sc_hd__conb_1 _332_ (
    .LO(io_out[5])
  );
  sky130_fd_sc_hd__conb_1 _333_ (
    .LO(io_out[7])
  );
  sky130_fd_sc_hd__conb_1 _334_ (
    .LO(io_out[8])
  );
  sky130_fd_sc_hd__conb_1 _335_ (
    .LO(io_out[9])
  );
  sky130_fd_sc_hd__conb_1 _336_ (
    .LO(io_out[10])
  );
  sky130_fd_sc_hd__conb_1 _337_ (
    .LO(io_out[11])
  );
  sky130_fd_sc_hd__conb_1 _338_ (
    .LO(io_out[12])
  );
  sky130_fd_sc_hd__conb_1 _339_ (
    .LO(io_out[14])
  );
  sky130_fd_sc_hd__conb_1 _340_ (
    .LO(io_out[27])
  );
  sky130_fd_sc_hd__conb_1 _341_ (
    .LO(io_out[28])
  );
  sky130_fd_sc_hd__conb_1 _342_ (
    .LO(io_out[29])
  );
  sky130_fd_sc_hd__conb_1 _343_ (
    .LO(io_out[30])
  );
  sky130_fd_sc_hd__conb_1 _344_ (
    .LO(io_out[31])
  );
  sky130_fd_sc_hd__conb_1 _345_ (
    .LO(io_out[32])
  );
  sky130_fd_sc_hd__conb_1 _346_ (
    .LO(io_out[33])
  );
  sky130_fd_sc_hd__conb_1 _347_ (
    .LO(io_out[34])
  );
  sky130_fd_sc_hd__conb_1 _348_ (
    .LO(io_out[35])
  );
  sky130_fd_sc_hd__conb_1 _349_ (
    .LO(io_out[36])
  );
  sky130_fd_sc_hd__conb_1 _350_ (
    .LO(io_out[37])
  );
  sky130_fd_sc_hd__buf_2 _351_ (
    .A(ReceiveLED),
    .X(io_out[6])
  );
  sky130_fd_sc_hd__buf_2 _352_ (
    .A(ComActive),
    .X(la_data_out[0])
  );
  sky130_fd_sc_hd__buf_2 _353_ (
    .A(io_in[5]),
    .X(la_data_out[1])
  );
  sky130_fd_sc_hd__buf_2 _354_ (
    .A(ReceiveLED),
    .X(la_data_out[2])
  );
  sky130_fd_sc_hd__mux2_1 _355_ (
    .A0(wb_clk_i),
    .A1(user_clock2),
    .S(io_in[2]),
    .X(_000_)
  );
  sky130_fd_sc_hd__mux2_1 _356_ (
    .A0(io_in[0]),
    .A1(_000_),
    .S(io_in[1]),
    .X(CLK)
  );
  sky130_fd_sc_hd__mux2_1 _357_ (
    .A0(la_data_in[0]),
    .A1(io_in[8]),
    .S(io_in[7]),
    .X(debug_req_1)
  );
  sky130_fd_sc_hd__mux2_1 _358_ (
    .A0(la_data_in[1]),
    .A1(io_in[9]),
    .S(io_in[7]),
    .X(fetch_enable_1)
  );
  sky130_fd_sc_hd__mux2_1 _359_ (
    .A0(la_data_in[2]),
    .A1(io_in[10]),
    .S(io_in[7]),
    .X(debug_req_2)
  );
  sky130_fd_sc_hd__mux2_1 _360_ (
    .A0(la_data_in[3]),
    .A1(io_in[11]),
    .S(io_in[7]),
    .X(fetch_enable_2)
  );
  Config Config_inst (
    .CLK(CLK),
    .ComActive(ComActive),
    .ConfigWriteData({ \LocalWriteData[31] , \LocalWriteData[30] , \LocalWriteData[29] , \LocalWriteData[28] , \LocalWriteData[27] , \LocalWriteData[26] , \LocalWriteData[25] , \LocalWriteData[24] , \LocalWriteData[23] , \LocalWriteData[22] , \LocalWriteData[21] , \LocalWriteData[20] , \LocalWriteData[19] , \LocalWriteData[18] , \LocalWriteData[17] , \LocalWriteData[16] , \LocalWriteData[15] , \LocalWriteData[14] , \LocalWriteData[13] , \LocalWriteData[12] , \LocalWriteData[11] , \LocalWriteData[10] , \LocalWriteData[9] , \LocalWriteData[8] , \LocalWriteData[7] , \LocalWriteData[6] , \LocalWriteData[5] , \LocalWriteData[4] , \LocalWriteData[3] , \LocalWriteData[2] , \LocalWriteData[1] , \LocalWriteData[0]  }),
    .ConfigWriteStrobe(LocalWriteStrobe),
    .FrameAddressRegister({ \FrameAddressRegister[31] , \FrameAddressRegister[30] , \FrameAddressRegister[29] , \FrameAddressRegister[28] , \FrameAddressRegister[27] , \FrameAddressRegister[26] , \FrameAddressRegister[25] , \FrameAddressRegister[24] , \FrameAddressRegister[23] , \FrameAddressRegister[22] , \FrameAddressRegister[21] , \FrameAddressRegister[20] , \FrameAddressRegister[19] , \FrameAddressRegister[18] , \FrameAddressRegister[17] , \FrameAddressRegister[16] , \FrameAddressRegister[15] , \FrameAddressRegister[14] , \FrameAddressRegister[13] , \FrameAddressRegister[12] , \FrameAddressRegister[11] , \FrameAddressRegister[10] , \FrameAddressRegister[9] , \FrameAddressRegister[8] , \FrameAddressRegister[7] , \FrameAddressRegister[6] , \FrameAddressRegister[5] , \FrameAddressRegister[4] , \FrameAddressRegister[3] , \FrameAddressRegister[2] , \FrameAddressRegister[1] , \FrameAddressRegister[0]  }),
    .LongFrameStrobe(LongFrameStrobe),
    .ReceiveLED(ReceiveLED),
    .RowSelect({ \RowSelect[4] , \RowSelect[3] , \RowSelect[2] , \RowSelect[1] , \RowSelect[0]  }),
    .Rx(io_in[5]),
    .SelfWriteData({ \SelfWriteData[31] , \SelfWriteData[30] , \SelfWriteData[29] , \SelfWriteData[28] , \SelfWriteData[27] , \SelfWriteData[26] , \SelfWriteData[25] , \SelfWriteData[24] , \SelfWriteData[23] , \SelfWriteData[22] , \SelfWriteData[21] , \SelfWriteData[20] , \SelfWriteData[19] , \SelfWriteData[18] , \SelfWriteData[17] , \SelfWriteData[16] , \SelfWriteData[15] , \SelfWriteData[14] , \SelfWriteData[13] , \SelfWriteData[12] , \SelfWriteData[11] , \SelfWriteData[10] , \SelfWriteData[9] , \SelfWriteData[8] , \SelfWriteData[7] , \SelfWriteData[6] , \SelfWriteData[5] , \SelfWriteData[4] , \SelfWriteData[3] , \SelfWriteData[2] , \SelfWriteData[1] , \SelfWriteData[0]  }),
    .SelfWriteStrobe(SelfWriteStrobe),
    .s_clk(io_in[3]),
    .s_data(io_in[4])
  );
  Frame_Data_Reg_0 Inst_Frame_Data_Reg_0 (
    .CLK(CLK),
    .FrameData_I({ \LocalWriteData[31] , \LocalWriteData[30] , \LocalWriteData[29] , \LocalWriteData[28] , \LocalWriteData[27] , \LocalWriteData[26] , \LocalWriteData[25] , \LocalWriteData[24] , \LocalWriteData[23] , \LocalWriteData[22] , \LocalWriteData[21] , \LocalWriteData[20] , \LocalWriteData[19] , \LocalWriteData[18] , \LocalWriteData[17] , \LocalWriteData[16] , \LocalWriteData[15] , \LocalWriteData[14] , \LocalWriteData[13] , \LocalWriteData[12] , \LocalWriteData[11] , \LocalWriteData[10] , \LocalWriteData[9] , \LocalWriteData[8] , \LocalWriteData[7] , \LocalWriteData[6] , \LocalWriteData[5] , \LocalWriteData[4] , \LocalWriteData[3] , \LocalWriteData[2] , \LocalWriteData[1] , \LocalWriteData[0]  }),
    .FrameData_O({ \FrameData[63] , \FrameData[62] , \FrameData[61] , \FrameData[60] , \FrameData[59] , \FrameData[58] , \FrameData[57] , \FrameData[56] , \FrameData[55] , \FrameData[54] , \FrameData[53] , \FrameData[52] , \FrameData[51] , \FrameData[50] , \FrameData[49] , \FrameData[48] , \FrameData[47] , \FrameData[46] , \FrameData[45] , \FrameData[44] , \FrameData[43] , \FrameData[42] , \FrameData[41] , \FrameData[40] , \FrameData[39] , \FrameData[38] , \FrameData[37] , \FrameData[36] , \FrameData[35] , \FrameData[34] , \FrameData[33] , \FrameData[32]  }),
    .RowSelect({ \RowSelect[4] , \RowSelect[3] , \RowSelect[2] , \RowSelect[1] , \RowSelect[0]  })
  );
  Frame_Data_Reg_1 Inst_Frame_Data_Reg_1 (
    .CLK(CLK),
    .FrameData_I({ \LocalWriteData[31] , \LocalWriteData[30] , \LocalWriteData[29] , \LocalWriteData[28] , \LocalWriteData[27] , \LocalWriteData[26] , \LocalWriteData[25] , \LocalWriteData[24] , \LocalWriteData[23] , \LocalWriteData[22] , \LocalWriteData[21] , \LocalWriteData[20] , \LocalWriteData[19] , \LocalWriteData[18] , \LocalWriteData[17] , \LocalWriteData[16] , \LocalWriteData[15] , \LocalWriteData[14] , \LocalWriteData[13] , \LocalWriteData[12] , \LocalWriteData[11] , \LocalWriteData[10] , \LocalWriteData[9] , \LocalWriteData[8] , \LocalWriteData[7] , \LocalWriteData[6] , \LocalWriteData[5] , \LocalWriteData[4] , \LocalWriteData[3] , \LocalWriteData[2] , \LocalWriteData[1] , \LocalWriteData[0]  }),
    .FrameData_O({ \FrameData[95] , \FrameData[94] , \FrameData[93] , \FrameData[92] , \FrameData[91] , \FrameData[90] , \FrameData[89] , \FrameData[88] , \FrameData[87] , \FrameData[86] , \FrameData[85] , \FrameData[84] , \FrameData[83] , \FrameData[82] , \FrameData[81] , \FrameData[80] , \FrameData[79] , \FrameData[78] , \FrameData[77] , \FrameData[76] , \FrameData[75] , \FrameData[74] , \FrameData[73] , \FrameData[72] , \FrameData[71] , \FrameData[70] , \FrameData[69] , \FrameData[68] , \FrameData[67] , \FrameData[66] , \FrameData[65] , \FrameData[64]  }),
    .RowSelect({ \RowSelect[4] , \RowSelect[3] , \RowSelect[2] , \RowSelect[1] , \RowSelect[0]  })
  );
  Frame_Data_Reg_10 Inst_Frame_Data_Reg_10 (
    .CLK(CLK),
    .FrameData_I({ \LocalWriteData[31] , \LocalWriteData[30] , \LocalWriteData[29] , \LocalWriteData[28] , \LocalWriteData[27] , \LocalWriteData[26] , \LocalWriteData[25] , \LocalWriteData[24] , \LocalWriteData[23] , \LocalWriteData[22] , \LocalWriteData[21] , \LocalWriteData[20] , \LocalWriteData[19] , \LocalWriteData[18] , \LocalWriteData[17] , \LocalWriteData[16] , \LocalWriteData[15] , \LocalWriteData[14] , \LocalWriteData[13] , \LocalWriteData[12] , \LocalWriteData[11] , \LocalWriteData[10] , \LocalWriteData[9] , \LocalWriteData[8] , \LocalWriteData[7] , \LocalWriteData[6] , \LocalWriteData[5] , \LocalWriteData[4] , \LocalWriteData[3] , \LocalWriteData[2] , \LocalWriteData[1] , \LocalWriteData[0]  }),
    .FrameData_O({ \FrameData[383] , \FrameData[382] , \FrameData[381] , \FrameData[380] , \FrameData[379] , \FrameData[378] , \FrameData[377] , \FrameData[376] , \FrameData[375] , \FrameData[374] , \FrameData[373] , \FrameData[372] , \FrameData[371] , \FrameData[370] , \FrameData[369] , \FrameData[368] , \FrameData[367] , \FrameData[366] , \FrameData[365] , \FrameData[364] , \FrameData[363] , \FrameData[362] , \FrameData[361] , \FrameData[360] , \FrameData[359] , \FrameData[358] , \FrameData[357] , \FrameData[356] , \FrameData[355] , \FrameData[354] , \FrameData[353] , \FrameData[352]  }),
    .RowSelect({ \RowSelect[4] , \RowSelect[3] , \RowSelect[2] , \RowSelect[1] , \RowSelect[0]  })
  );
  Frame_Data_Reg_11 Inst_Frame_Data_Reg_11 (
    .CLK(CLK),
    .FrameData_I({ \LocalWriteData[31] , \LocalWriteData[30] , \LocalWriteData[29] , \LocalWriteData[28] , \LocalWriteData[27] , \LocalWriteData[26] , \LocalWriteData[25] , \LocalWriteData[24] , \LocalWriteData[23] , \LocalWriteData[22] , \LocalWriteData[21] , \LocalWriteData[20] , \LocalWriteData[19] , \LocalWriteData[18] , \LocalWriteData[17] , \LocalWriteData[16] , \LocalWriteData[15] , \LocalWriteData[14] , \LocalWriteData[13] , \LocalWriteData[12] , \LocalWriteData[11] , \LocalWriteData[10] , \LocalWriteData[9] , \LocalWriteData[8] , \LocalWriteData[7] , \LocalWriteData[6] , \LocalWriteData[5] , \LocalWriteData[4] , \LocalWriteData[3] , \LocalWriteData[2] , \LocalWriteData[1] , \LocalWriteData[0]  }),
    .FrameData_O({ \FrameData[415] , \FrameData[414] , \FrameData[413] , \FrameData[412] , \FrameData[411] , \FrameData[410] , \FrameData[409] , \FrameData[408] , \FrameData[407] , \FrameData[406] , \FrameData[405] , \FrameData[404] , \FrameData[403] , \FrameData[402] , \FrameData[401] , \FrameData[400] , \FrameData[399] , \FrameData[398] , \FrameData[397] , \FrameData[396] , \FrameData[395] , \FrameData[394] , \FrameData[393] , \FrameData[392] , \FrameData[391] , \FrameData[390] , \FrameData[389] , \FrameData[388] , \FrameData[387] , \FrameData[386] , \FrameData[385] , \FrameData[384]  }),
    .RowSelect({ \RowSelect[4] , \RowSelect[3] , \RowSelect[2] , \RowSelect[1] , \RowSelect[0]  })
  );
  Frame_Data_Reg_12 Inst_Frame_Data_Reg_12 (
    .CLK(CLK),
    .FrameData_I({ \LocalWriteData[31] , \LocalWriteData[30] , \LocalWriteData[29] , \LocalWriteData[28] , \LocalWriteData[27] , \LocalWriteData[26] , \LocalWriteData[25] , \LocalWriteData[24] , \LocalWriteData[23] , \LocalWriteData[22] , \LocalWriteData[21] , \LocalWriteData[20] , \LocalWriteData[19] , \LocalWriteData[18] , \LocalWriteData[17] , \LocalWriteData[16] , \LocalWriteData[15] , \LocalWriteData[14] , \LocalWriteData[13] , \LocalWriteData[12] , \LocalWriteData[11] , \LocalWriteData[10] , \LocalWriteData[9] , \LocalWriteData[8] , \LocalWriteData[7] , \LocalWriteData[6] , \LocalWriteData[5] , \LocalWriteData[4] , \LocalWriteData[3] , \LocalWriteData[2] , \LocalWriteData[1] , \LocalWriteData[0]  }),
    .FrameData_O({ \FrameData[447] , \FrameData[446] , \FrameData[445] , \FrameData[444] , \FrameData[443] , \FrameData[442] , \FrameData[441] , \FrameData[440] , \FrameData[439] , \FrameData[438] , \FrameData[437] , \FrameData[436] , \FrameData[435] , \FrameData[434] , \FrameData[433] , \FrameData[432] , \FrameData[431] , \FrameData[430] , \FrameData[429] , \FrameData[428] , \FrameData[427] , \FrameData[426] , \FrameData[425] , \FrameData[424] , \FrameData[423] , \FrameData[422] , \FrameData[421] , \FrameData[420] , \FrameData[419] , \FrameData[418] , \FrameData[417] , \FrameData[416]  }),
    .RowSelect({ \RowSelect[4] , \RowSelect[3] , \RowSelect[2] , \RowSelect[1] , \RowSelect[0]  })
  );
  Frame_Data_Reg_13 Inst_Frame_Data_Reg_13 (
    .CLK(CLK),
    .FrameData_I({ \LocalWriteData[31] , \LocalWriteData[30] , \LocalWriteData[29] , \LocalWriteData[28] , \LocalWriteData[27] , \LocalWriteData[26] , \LocalWriteData[25] , \LocalWriteData[24] , \LocalWriteData[23] , \LocalWriteData[22] , \LocalWriteData[21] , \LocalWriteData[20] , \LocalWriteData[19] , \LocalWriteData[18] , \LocalWriteData[17] , \LocalWriteData[16] , \LocalWriteData[15] , \LocalWriteData[14] , \LocalWriteData[13] , \LocalWriteData[12] , \LocalWriteData[11] , \LocalWriteData[10] , \LocalWriteData[9] , \LocalWriteData[8] , \LocalWriteData[7] , \LocalWriteData[6] , \LocalWriteData[5] , \LocalWriteData[4] , \LocalWriteData[3] , \LocalWriteData[2] , \LocalWriteData[1] , \LocalWriteData[0]  }),
    .FrameData_O({ \FrameData[479] , \FrameData[478] , \FrameData[477] , \FrameData[476] , \FrameData[475] , \FrameData[474] , \FrameData[473] , \FrameData[472] , \FrameData[471] , \FrameData[470] , \FrameData[469] , \FrameData[468] , \FrameData[467] , \FrameData[466] , \FrameData[465] , \FrameData[464] , \FrameData[463] , \FrameData[462] , \FrameData[461] , \FrameData[460] , \FrameData[459] , \FrameData[458] , \FrameData[457] , \FrameData[456] , \FrameData[455] , \FrameData[454] , \FrameData[453] , \FrameData[452] , \FrameData[451] , \FrameData[450] , \FrameData[449] , \FrameData[448]  }),
    .RowSelect({ \RowSelect[4] , \RowSelect[3] , \RowSelect[2] , \RowSelect[1] , \RowSelect[0]  })
  );
  Frame_Data_Reg_2 Inst_Frame_Data_Reg_2 (
    .CLK(CLK),
    .FrameData_I({ \LocalWriteData[31] , \LocalWriteData[30] , \LocalWriteData[29] , \LocalWriteData[28] , \LocalWriteData[27] , \LocalWriteData[26] , \LocalWriteData[25] , \LocalWriteData[24] , \LocalWriteData[23] , \LocalWriteData[22] , \LocalWriteData[21] , \LocalWriteData[20] , \LocalWriteData[19] , \LocalWriteData[18] , \LocalWriteData[17] , \LocalWriteData[16] , \LocalWriteData[15] , \LocalWriteData[14] , \LocalWriteData[13] , \LocalWriteData[12] , \LocalWriteData[11] , \LocalWriteData[10] , \LocalWriteData[9] , \LocalWriteData[8] , \LocalWriteData[7] , \LocalWriteData[6] , \LocalWriteData[5] , \LocalWriteData[4] , \LocalWriteData[3] , \LocalWriteData[2] , \LocalWriteData[1] , \LocalWriteData[0]  }),
    .FrameData_O({ \FrameData[127] , \FrameData[126] , \FrameData[125] , \FrameData[124] , \FrameData[123] , \FrameData[122] , \FrameData[121] , \FrameData[120] , \FrameData[119] , \FrameData[118] , \FrameData[117] , \FrameData[116] , \FrameData[115] , \FrameData[114] , \FrameData[113] , \FrameData[112] , \FrameData[111] , \FrameData[110] , \FrameData[109] , \FrameData[108] , \FrameData[107] , \FrameData[106] , \FrameData[105] , \FrameData[104] , \FrameData[103] , \FrameData[102] , \FrameData[101] , \FrameData[100] , \FrameData[99] , \FrameData[98] , \FrameData[97] , \FrameData[96]  }),
    .RowSelect({ \RowSelect[4] , \RowSelect[3] , \RowSelect[2] , \RowSelect[1] , \RowSelect[0]  })
  );
  Frame_Data_Reg_3 Inst_Frame_Data_Reg_3 (
    .CLK(CLK),
    .FrameData_I({ \LocalWriteData[31] , \LocalWriteData[30] , \LocalWriteData[29] , \LocalWriteData[28] , \LocalWriteData[27] , \LocalWriteData[26] , \LocalWriteData[25] , \LocalWriteData[24] , \LocalWriteData[23] , \LocalWriteData[22] , \LocalWriteData[21] , \LocalWriteData[20] , \LocalWriteData[19] , \LocalWriteData[18] , \LocalWriteData[17] , \LocalWriteData[16] , \LocalWriteData[15] , \LocalWriteData[14] , \LocalWriteData[13] , \LocalWriteData[12] , \LocalWriteData[11] , \LocalWriteData[10] , \LocalWriteData[9] , \LocalWriteData[8] , \LocalWriteData[7] , \LocalWriteData[6] , \LocalWriteData[5] , \LocalWriteData[4] , \LocalWriteData[3] , \LocalWriteData[2] , \LocalWriteData[1] , \LocalWriteData[0]  }),
    .FrameData_O({ \FrameData[159] , \FrameData[158] , \FrameData[157] , \FrameData[156] , \FrameData[155] , \FrameData[154] , \FrameData[153] , \FrameData[152] , \FrameData[151] , \FrameData[150] , \FrameData[149] , \FrameData[148] , \FrameData[147] , \FrameData[146] , \FrameData[145] , \FrameData[144] , \FrameData[143] , \FrameData[142] , \FrameData[141] , \FrameData[140] , \FrameData[139] , \FrameData[138] , \FrameData[137] , \FrameData[136] , \FrameData[135] , \FrameData[134] , \FrameData[133] , \FrameData[132] , \FrameData[131] , \FrameData[130] , \FrameData[129] , \FrameData[128]  }),
    .RowSelect({ \RowSelect[4] , \RowSelect[3] , \RowSelect[2] , \RowSelect[1] , \RowSelect[0]  })
  );
  Frame_Data_Reg_4 Inst_Frame_Data_Reg_4 (
    .CLK(CLK),
    .FrameData_I({ \LocalWriteData[31] , \LocalWriteData[30] , \LocalWriteData[29] , \LocalWriteData[28] , \LocalWriteData[27] , \LocalWriteData[26] , \LocalWriteData[25] , \LocalWriteData[24] , \LocalWriteData[23] , \LocalWriteData[22] , \LocalWriteData[21] , \LocalWriteData[20] , \LocalWriteData[19] , \LocalWriteData[18] , \LocalWriteData[17] , \LocalWriteData[16] , \LocalWriteData[15] , \LocalWriteData[14] , \LocalWriteData[13] , \LocalWriteData[12] , \LocalWriteData[11] , \LocalWriteData[10] , \LocalWriteData[9] , \LocalWriteData[8] , \LocalWriteData[7] , \LocalWriteData[6] , \LocalWriteData[5] , \LocalWriteData[4] , \LocalWriteData[3] , \LocalWriteData[2] , \LocalWriteData[1] , \LocalWriteData[0]  }),
    .FrameData_O({ \FrameData[191] , \FrameData[190] , \FrameData[189] , \FrameData[188] , \FrameData[187] , \FrameData[186] , \FrameData[185] , \FrameData[184] , \FrameData[183] , \FrameData[182] , \FrameData[181] , \FrameData[180] , \FrameData[179] , \FrameData[178] , \FrameData[177] , \FrameData[176] , \FrameData[175] , \FrameData[174] , \FrameData[173] , \FrameData[172] , \FrameData[171] , \FrameData[170] , \FrameData[169] , \FrameData[168] , \FrameData[167] , \FrameData[166] , \FrameData[165] , \FrameData[164] , \FrameData[163] , \FrameData[162] , \FrameData[161] , \FrameData[160]  }),
    .RowSelect({ \RowSelect[4] , \RowSelect[3] , \RowSelect[2] , \RowSelect[1] , \RowSelect[0]  })
  );
  Frame_Data_Reg_5 Inst_Frame_Data_Reg_5 (
    .CLK(CLK),
    .FrameData_I({ \LocalWriteData[31] , \LocalWriteData[30] , \LocalWriteData[29] , \LocalWriteData[28] , \LocalWriteData[27] , \LocalWriteData[26] , \LocalWriteData[25] , \LocalWriteData[24] , \LocalWriteData[23] , \LocalWriteData[22] , \LocalWriteData[21] , \LocalWriteData[20] , \LocalWriteData[19] , \LocalWriteData[18] , \LocalWriteData[17] , \LocalWriteData[16] , \LocalWriteData[15] , \LocalWriteData[14] , \LocalWriteData[13] , \LocalWriteData[12] , \LocalWriteData[11] , \LocalWriteData[10] , \LocalWriteData[9] , \LocalWriteData[8] , \LocalWriteData[7] , \LocalWriteData[6] , \LocalWriteData[5] , \LocalWriteData[4] , \LocalWriteData[3] , \LocalWriteData[2] , \LocalWriteData[1] , \LocalWriteData[0]  }),
    .FrameData_O({ \FrameData[223] , \FrameData[222] , \FrameData[221] , \FrameData[220] , \FrameData[219] , \FrameData[218] , \FrameData[217] , \FrameData[216] , \FrameData[215] , \FrameData[214] , \FrameData[213] , \FrameData[212] , \FrameData[211] , \FrameData[210] , \FrameData[209] , \FrameData[208] , \FrameData[207] , \FrameData[206] , \FrameData[205] , \FrameData[204] , \FrameData[203] , \FrameData[202] , \FrameData[201] , \FrameData[200] , \FrameData[199] , \FrameData[198] , \FrameData[197] , \FrameData[196] , \FrameData[195] , \FrameData[194] , \FrameData[193] , \FrameData[192]  }),
    .RowSelect({ \RowSelect[4] , \RowSelect[3] , \RowSelect[2] , \RowSelect[1] , \RowSelect[0]  })
  );
  Frame_Data_Reg_6 Inst_Frame_Data_Reg_6 (
    .CLK(CLK),
    .FrameData_I({ \LocalWriteData[31] , \LocalWriteData[30] , \LocalWriteData[29] , \LocalWriteData[28] , \LocalWriteData[27] , \LocalWriteData[26] , \LocalWriteData[25] , \LocalWriteData[24] , \LocalWriteData[23] , \LocalWriteData[22] , \LocalWriteData[21] , \LocalWriteData[20] , \LocalWriteData[19] , \LocalWriteData[18] , \LocalWriteData[17] , \LocalWriteData[16] , \LocalWriteData[15] , \LocalWriteData[14] , \LocalWriteData[13] , \LocalWriteData[12] , \LocalWriteData[11] , \LocalWriteData[10] , \LocalWriteData[9] , \LocalWriteData[8] , \LocalWriteData[7] , \LocalWriteData[6] , \LocalWriteData[5] , \LocalWriteData[4] , \LocalWriteData[3] , \LocalWriteData[2] , \LocalWriteData[1] , \LocalWriteData[0]  }),
    .FrameData_O({ \FrameData[255] , \FrameData[254] , \FrameData[253] , \FrameData[252] , \FrameData[251] , \FrameData[250] , \FrameData[249] , \FrameData[248] , \FrameData[247] , \FrameData[246] , \FrameData[245] , \FrameData[244] , \FrameData[243] , \FrameData[242] , \FrameData[241] , \FrameData[240] , \FrameData[239] , \FrameData[238] , \FrameData[237] , \FrameData[236] , \FrameData[235] , \FrameData[234] , \FrameData[233] , \FrameData[232] , \FrameData[231] , \FrameData[230] , \FrameData[229] , \FrameData[228] , \FrameData[227] , \FrameData[226] , \FrameData[225] , \FrameData[224]  }),
    .RowSelect({ \RowSelect[4] , \RowSelect[3] , \RowSelect[2] , \RowSelect[1] , \RowSelect[0]  })
  );
  Frame_Data_Reg_7 Inst_Frame_Data_Reg_7 (
    .CLK(CLK),
    .FrameData_I({ \LocalWriteData[31] , \LocalWriteData[30] , \LocalWriteData[29] , \LocalWriteData[28] , \LocalWriteData[27] , \LocalWriteData[26] , \LocalWriteData[25] , \LocalWriteData[24] , \LocalWriteData[23] , \LocalWriteData[22] , \LocalWriteData[21] , \LocalWriteData[20] , \LocalWriteData[19] , \LocalWriteData[18] , \LocalWriteData[17] , \LocalWriteData[16] , \LocalWriteData[15] , \LocalWriteData[14] , \LocalWriteData[13] , \LocalWriteData[12] , \LocalWriteData[11] , \LocalWriteData[10] , \LocalWriteData[9] , \LocalWriteData[8] , \LocalWriteData[7] , \LocalWriteData[6] , \LocalWriteData[5] , \LocalWriteData[4] , \LocalWriteData[3] , \LocalWriteData[2] , \LocalWriteData[1] , \LocalWriteData[0]  }),
    .FrameData_O({ \FrameData[287] , \FrameData[286] , \FrameData[285] , \FrameData[284] , \FrameData[283] , \FrameData[282] , \FrameData[281] , \FrameData[280] , \FrameData[279] , \FrameData[278] , \FrameData[277] , \FrameData[276] , \FrameData[275] , \FrameData[274] , \FrameData[273] , \FrameData[272] , \FrameData[271] , \FrameData[270] , \FrameData[269] , \FrameData[268] , \FrameData[267] , \FrameData[266] , \FrameData[265] , \FrameData[264] , \FrameData[263] , \FrameData[262] , \FrameData[261] , \FrameData[260] , \FrameData[259] , \FrameData[258] , \FrameData[257] , \FrameData[256]  }),
    .RowSelect({ \RowSelect[4] , \RowSelect[3] , \RowSelect[2] , \RowSelect[1] , \RowSelect[0]  })
  );
  Frame_Data_Reg_8 Inst_Frame_Data_Reg_8 (
    .CLK(CLK),
    .FrameData_I({ \LocalWriteData[31] , \LocalWriteData[30] , \LocalWriteData[29] , \LocalWriteData[28] , \LocalWriteData[27] , \LocalWriteData[26] , \LocalWriteData[25] , \LocalWriteData[24] , \LocalWriteData[23] , \LocalWriteData[22] , \LocalWriteData[21] , \LocalWriteData[20] , \LocalWriteData[19] , \LocalWriteData[18] , \LocalWriteData[17] , \LocalWriteData[16] , \LocalWriteData[15] , \LocalWriteData[14] , \LocalWriteData[13] , \LocalWriteData[12] , \LocalWriteData[11] , \LocalWriteData[10] , \LocalWriteData[9] , \LocalWriteData[8] , \LocalWriteData[7] , \LocalWriteData[6] , \LocalWriteData[5] , \LocalWriteData[4] , \LocalWriteData[3] , \LocalWriteData[2] , \LocalWriteData[1] , \LocalWriteData[0]  }),
    .FrameData_O({ \FrameData[319] , \FrameData[318] , \FrameData[317] , \FrameData[316] , \FrameData[315] , \FrameData[314] , \FrameData[313] , \FrameData[312] , \FrameData[311] , \FrameData[310] , \FrameData[309] , \FrameData[308] , \FrameData[307] , \FrameData[306] , \FrameData[305] , \FrameData[304] , \FrameData[303] , \FrameData[302] , \FrameData[301] , \FrameData[300] , \FrameData[299] , \FrameData[298] , \FrameData[297] , \FrameData[296] , \FrameData[295] , \FrameData[294] , \FrameData[293] , \FrameData[292] , \FrameData[291] , \FrameData[290] , \FrameData[289] , \FrameData[288]  }),
    .RowSelect({ \RowSelect[4] , \RowSelect[3] , \RowSelect[2] , \RowSelect[1] , \RowSelect[0]  })
  );
  Frame_Data_Reg_9 Inst_Frame_Data_Reg_9 (
    .CLK(CLK),
    .FrameData_I({ \LocalWriteData[31] , \LocalWriteData[30] , \LocalWriteData[29] , \LocalWriteData[28] , \LocalWriteData[27] , \LocalWriteData[26] , \LocalWriteData[25] , \LocalWriteData[24] , \LocalWriteData[23] , \LocalWriteData[22] , \LocalWriteData[21] , \LocalWriteData[20] , \LocalWriteData[19] , \LocalWriteData[18] , \LocalWriteData[17] , \LocalWriteData[16] , \LocalWriteData[15] , \LocalWriteData[14] , \LocalWriteData[13] , \LocalWriteData[12] , \LocalWriteData[11] , \LocalWriteData[10] , \LocalWriteData[9] , \LocalWriteData[8] , \LocalWriteData[7] , \LocalWriteData[6] , \LocalWriteData[5] , \LocalWriteData[4] , \LocalWriteData[3] , \LocalWriteData[2] , \LocalWriteData[1] , \LocalWriteData[0]  }),
    .FrameData_O({ \FrameData[351] , \FrameData[350] , \FrameData[349] , \FrameData[348] , \FrameData[347] , \FrameData[346] , \FrameData[345] , \FrameData[344] , \FrameData[343] , \FrameData[342] , \FrameData[341] , \FrameData[340] , \FrameData[339] , \FrameData[338] , \FrameData[337] , \FrameData[336] , \FrameData[335] , \FrameData[334] , \FrameData[333] , \FrameData[332] , \FrameData[331] , \FrameData[330] , \FrameData[329] , \FrameData[328] , \FrameData[327] , \FrameData[326] , \FrameData[325] , \FrameData[324] , \FrameData[323] , \FrameData[322] , \FrameData[321] , \FrameData[320]  }),
    .RowSelect({ \RowSelect[4] , \RowSelect[3] , \RowSelect[2] , \RowSelect[1] , \RowSelect[0]  })
  );
  Frame_Select_0 Inst_Frame_Select_0 (
    .FrameSelect({ \FrameAddressRegister[31] , \FrameAddressRegister[30] , \FrameAddressRegister[29] , \FrameAddressRegister[28] , \FrameAddressRegister[27]  }),
    .FrameStrobe(LongFrameStrobe),
    .FrameStrobe_I({ \FrameAddressRegister[19] , \FrameAddressRegister[18] , \FrameAddressRegister[17] , \FrameAddressRegister[16] , \FrameAddressRegister[15] , \FrameAddressRegister[14] , \FrameAddressRegister[13] , \FrameAddressRegister[12] , \FrameAddressRegister[11] , \FrameAddressRegister[10] , \FrameAddressRegister[9] , \FrameAddressRegister[8] , \FrameAddressRegister[7] , \FrameAddressRegister[6] , \FrameAddressRegister[5] , \FrameAddressRegister[4] , \FrameAddressRegister[3] , \FrameAddressRegister[2] , \FrameAddressRegister[1] , \FrameAddressRegister[0]  }),
    .FrameStrobe_O({ \FrameSelect[19] , \FrameSelect[18] , \FrameSelect[17] , \FrameSelect[16] , \FrameSelect[15] , \FrameSelect[14] , \FrameSelect[13] , \FrameSelect[12] , \FrameSelect[11] , \FrameSelect[10] , \FrameSelect[9] , \FrameSelect[8] , \FrameSelect[7] , \FrameSelect[6] , \FrameSelect[5] , \FrameSelect[4] , \FrameSelect[3] , \FrameSelect[2] , \FrameSelect[1] , \FrameSelect[0]  })
  );
  Frame_Select_1 Inst_Frame_Select_1 (
    .FrameSelect({ \FrameAddressRegister[31] , \FrameAddressRegister[30] , \FrameAddressRegister[29] , \FrameAddressRegister[28] , \FrameAddressRegister[27]  }),
    .FrameStrobe(LongFrameStrobe),
    .FrameStrobe_I({ \FrameAddressRegister[19] , \FrameAddressRegister[18] , \FrameAddressRegister[17] , \FrameAddressRegister[16] , \FrameAddressRegister[15] , \FrameAddressRegister[14] , \FrameAddressRegister[13] , \FrameAddressRegister[12] , \FrameAddressRegister[11] , \FrameAddressRegister[10] , \FrameAddressRegister[9] , \FrameAddressRegister[8] , \FrameAddressRegister[7] , \FrameAddressRegister[6] , \FrameAddressRegister[5] , \FrameAddressRegister[4] , \FrameAddressRegister[3] , \FrameAddressRegister[2] , \FrameAddressRegister[1] , \FrameAddressRegister[0]  }),
    .FrameStrobe_O({ \FrameSelect[39] , \FrameSelect[38] , \FrameSelect[37] , \FrameSelect[36] , \FrameSelect[35] , \FrameSelect[34] , \FrameSelect[33] , \FrameSelect[32] , \FrameSelect[31] , \FrameSelect[30] , \FrameSelect[29] , \FrameSelect[28] , \FrameSelect[27] , \FrameSelect[26] , \FrameSelect[25] , \FrameSelect[24] , \FrameSelect[23] , \FrameSelect[22] , \FrameSelect[21] , \FrameSelect[20]  })
  );
  Frame_Select_10 Inst_Frame_Select_10 (
    .FrameSelect({ \FrameAddressRegister[31] , \FrameAddressRegister[30] , \FrameAddressRegister[29] , \FrameAddressRegister[28] , \FrameAddressRegister[27]  }),
    .FrameStrobe(LongFrameStrobe),
    .FrameStrobe_I({ \FrameAddressRegister[19] , \FrameAddressRegister[18] , \FrameAddressRegister[17] , \FrameAddressRegister[16] , \FrameAddressRegister[15] , \FrameAddressRegister[14] , \FrameAddressRegister[13] , \FrameAddressRegister[12] , \FrameAddressRegister[11] , \FrameAddressRegister[10] , \FrameAddressRegister[9] , \FrameAddressRegister[8] , \FrameAddressRegister[7] , \FrameAddressRegister[6] , \FrameAddressRegister[5] , \FrameAddressRegister[4] , \FrameAddressRegister[3] , \FrameAddressRegister[2] , \FrameAddressRegister[1] , \FrameAddressRegister[0]  }),
    .FrameStrobe_O({ \FrameSelect[219] , \FrameSelect[218] , \FrameSelect[217] , \FrameSelect[216] , \FrameSelect[215] , \FrameSelect[214] , \FrameSelect[213] , \FrameSelect[212] , \FrameSelect[211] , \FrameSelect[210] , \FrameSelect[209] , \FrameSelect[208] , \FrameSelect[207] , \FrameSelect[206] , \FrameSelect[205] , \FrameSelect[204] , \FrameSelect[203] , \FrameSelect[202] , \FrameSelect[201] , \FrameSelect[200]  })
  );
  Frame_Select_11 Inst_Frame_Select_11 (
    .FrameSelect({ \FrameAddressRegister[31] , \FrameAddressRegister[30] , \FrameAddressRegister[29] , \FrameAddressRegister[28] , \FrameAddressRegister[27]  }),
    .FrameStrobe(LongFrameStrobe),
    .FrameStrobe_I({ \FrameAddressRegister[19] , \FrameAddressRegister[18] , \FrameAddressRegister[17] , \FrameAddressRegister[16] , \FrameAddressRegister[15] , \FrameAddressRegister[14] , \FrameAddressRegister[13] , \FrameAddressRegister[12] , \FrameAddressRegister[11] , \FrameAddressRegister[10] , \FrameAddressRegister[9] , \FrameAddressRegister[8] , \FrameAddressRegister[7] , \FrameAddressRegister[6] , \FrameAddressRegister[5] , \FrameAddressRegister[4] , \FrameAddressRegister[3] , \FrameAddressRegister[2] , \FrameAddressRegister[1] , \FrameAddressRegister[0]  }),
    .FrameStrobe_O({ \FrameSelect[239] , \FrameSelect[238] , \FrameSelect[237] , \FrameSelect[236] , \FrameSelect[235] , \FrameSelect[234] , \FrameSelect[233] , \FrameSelect[232] , \FrameSelect[231] , \FrameSelect[230] , \FrameSelect[229] , \FrameSelect[228] , \FrameSelect[227] , \FrameSelect[226] , \FrameSelect[225] , \FrameSelect[224] , \FrameSelect[223] , \FrameSelect[222] , \FrameSelect[221] , \FrameSelect[220]  })
  );
  Frame_Select_12 Inst_Frame_Select_12 (
    .FrameSelect({ \FrameAddressRegister[31] , \FrameAddressRegister[30] , \FrameAddressRegister[29] , \FrameAddressRegister[28] , \FrameAddressRegister[27]  }),
    .FrameStrobe(LongFrameStrobe),
    .FrameStrobe_I({ \FrameAddressRegister[19] , \FrameAddressRegister[18] , \FrameAddressRegister[17] , \FrameAddressRegister[16] , \FrameAddressRegister[15] , \FrameAddressRegister[14] , \FrameAddressRegister[13] , \FrameAddressRegister[12] , \FrameAddressRegister[11] , \FrameAddressRegister[10] , \FrameAddressRegister[9] , \FrameAddressRegister[8] , \FrameAddressRegister[7] , \FrameAddressRegister[6] , \FrameAddressRegister[5] , \FrameAddressRegister[4] , \FrameAddressRegister[3] , \FrameAddressRegister[2] , \FrameAddressRegister[1] , \FrameAddressRegister[0]  }),
    .FrameStrobe_O({ \FrameSelect[259] , \FrameSelect[258] , \FrameSelect[257] , \FrameSelect[256] , \FrameSelect[255] , \FrameSelect[254] , \FrameSelect[253] , \FrameSelect[252] , \FrameSelect[251] , \FrameSelect[250] , \FrameSelect[249] , \FrameSelect[248] , \FrameSelect[247] , \FrameSelect[246] , \FrameSelect[245] , \FrameSelect[244] , \FrameSelect[243] , \FrameSelect[242] , \FrameSelect[241] , \FrameSelect[240]  })
  );
  Frame_Select_13 Inst_Frame_Select_13 (
    .FrameSelect({ \FrameAddressRegister[31] , \FrameAddressRegister[30] , \FrameAddressRegister[29] , \FrameAddressRegister[28] , \FrameAddressRegister[27]  }),
    .FrameStrobe(LongFrameStrobe),
    .FrameStrobe_I({ \FrameAddressRegister[19] , \FrameAddressRegister[18] , \FrameAddressRegister[17] , \FrameAddressRegister[16] , \FrameAddressRegister[15] , \FrameAddressRegister[14] , \FrameAddressRegister[13] , \FrameAddressRegister[12] , \FrameAddressRegister[11] , \FrameAddressRegister[10] , \FrameAddressRegister[9] , \FrameAddressRegister[8] , \FrameAddressRegister[7] , \FrameAddressRegister[6] , \FrameAddressRegister[5] , \FrameAddressRegister[4] , \FrameAddressRegister[3] , \FrameAddressRegister[2] , \FrameAddressRegister[1] , \FrameAddressRegister[0]  }),
    .FrameStrobe_O({ \FrameSelect[279] , \FrameSelect[278] , \FrameSelect[277] , \FrameSelect[276] , \FrameSelect[275] , \FrameSelect[274] , \FrameSelect[273] , \FrameSelect[272] , \FrameSelect[271] , \FrameSelect[270] , \FrameSelect[269] , \FrameSelect[268] , \FrameSelect[267] , \FrameSelect[266] , \FrameSelect[265] , \FrameSelect[264] , \FrameSelect[263] , \FrameSelect[262] , \FrameSelect[261] , \FrameSelect[260]  })
  );
  Frame_Select_14 Inst_Frame_Select_14 (
    .FrameSelect({ \FrameAddressRegister[31] , \FrameAddressRegister[30] , \FrameAddressRegister[29] , \FrameAddressRegister[28] , \FrameAddressRegister[27]  }),
    .FrameStrobe(LongFrameStrobe),
    .FrameStrobe_I({ \FrameAddressRegister[19] , \FrameAddressRegister[18] , \FrameAddressRegister[17] , \FrameAddressRegister[16] , \FrameAddressRegister[15] , \FrameAddressRegister[14] , \FrameAddressRegister[13] , \FrameAddressRegister[12] , \FrameAddressRegister[11] , \FrameAddressRegister[10] , \FrameAddressRegister[9] , \FrameAddressRegister[8] , \FrameAddressRegister[7] , \FrameAddressRegister[6] , \FrameAddressRegister[5] , \FrameAddressRegister[4] , \FrameAddressRegister[3] , \FrameAddressRegister[2] , \FrameAddressRegister[1] , \FrameAddressRegister[0]  }),
    .FrameStrobe_O({ \FrameSelect[299] , \FrameSelect[298] , \FrameSelect[297] , \FrameSelect[296] , \FrameSelect[295] , \FrameSelect[294] , \FrameSelect[293] , \FrameSelect[292] , \FrameSelect[291] , \FrameSelect[290] , \FrameSelect[289] , \FrameSelect[288] , \FrameSelect[287] , \FrameSelect[286] , \FrameSelect[285] , \FrameSelect[284] , \FrameSelect[283] , \FrameSelect[282] , \FrameSelect[281] , \FrameSelect[280]  })
  );
  Frame_Select_2 Inst_Frame_Select_2 (
    .FrameSelect({ \FrameAddressRegister[31] , \FrameAddressRegister[30] , \FrameAddressRegister[29] , \FrameAddressRegister[28] , \FrameAddressRegister[27]  }),
    .FrameStrobe(LongFrameStrobe),
    .FrameStrobe_I({ \FrameAddressRegister[19] , \FrameAddressRegister[18] , \FrameAddressRegister[17] , \FrameAddressRegister[16] , \FrameAddressRegister[15] , \FrameAddressRegister[14] , \FrameAddressRegister[13] , \FrameAddressRegister[12] , \FrameAddressRegister[11] , \FrameAddressRegister[10] , \FrameAddressRegister[9] , \FrameAddressRegister[8] , \FrameAddressRegister[7] , \FrameAddressRegister[6] , \FrameAddressRegister[5] , \FrameAddressRegister[4] , \FrameAddressRegister[3] , \FrameAddressRegister[2] , \FrameAddressRegister[1] , \FrameAddressRegister[0]  }),
    .FrameStrobe_O({ \FrameSelect[59] , \FrameSelect[58] , \FrameSelect[57] , \FrameSelect[56] , \FrameSelect[55] , \FrameSelect[54] , \FrameSelect[53] , \FrameSelect[52] , \FrameSelect[51] , \FrameSelect[50] , \FrameSelect[49] , \FrameSelect[48] , \FrameSelect[47] , \FrameSelect[46] , \FrameSelect[45] , \FrameSelect[44] , \FrameSelect[43] , \FrameSelect[42] , \FrameSelect[41] , \FrameSelect[40]  })
  );
  Frame_Select_3 Inst_Frame_Select_3 (
    .FrameSelect({ \FrameAddressRegister[31] , \FrameAddressRegister[30] , \FrameAddressRegister[29] , \FrameAddressRegister[28] , \FrameAddressRegister[27]  }),
    .FrameStrobe(LongFrameStrobe),
    .FrameStrobe_I({ \FrameAddressRegister[19] , \FrameAddressRegister[18] , \FrameAddressRegister[17] , \FrameAddressRegister[16] , \FrameAddressRegister[15] , \FrameAddressRegister[14] , \FrameAddressRegister[13] , \FrameAddressRegister[12] , \FrameAddressRegister[11] , \FrameAddressRegister[10] , \FrameAddressRegister[9] , \FrameAddressRegister[8] , \FrameAddressRegister[7] , \FrameAddressRegister[6] , \FrameAddressRegister[5] , \FrameAddressRegister[4] , \FrameAddressRegister[3] , \FrameAddressRegister[2] , \FrameAddressRegister[1] , \FrameAddressRegister[0]  }),
    .FrameStrobe_O({ \FrameSelect[79] , \FrameSelect[78] , \FrameSelect[77] , \FrameSelect[76] , \FrameSelect[75] , \FrameSelect[74] , \FrameSelect[73] , \FrameSelect[72] , \FrameSelect[71] , \FrameSelect[70] , \FrameSelect[69] , \FrameSelect[68] , \FrameSelect[67] , \FrameSelect[66] , \FrameSelect[65] , \FrameSelect[64] , \FrameSelect[63] , \FrameSelect[62] , \FrameSelect[61] , \FrameSelect[60]  })
  );
  Frame_Select_4 Inst_Frame_Select_4 (
    .FrameSelect({ \FrameAddressRegister[31] , \FrameAddressRegister[30] , \FrameAddressRegister[29] , \FrameAddressRegister[28] , \FrameAddressRegister[27]  }),
    .FrameStrobe(LongFrameStrobe),
    .FrameStrobe_I({ \FrameAddressRegister[19] , \FrameAddressRegister[18] , \FrameAddressRegister[17] , \FrameAddressRegister[16] , \FrameAddressRegister[15] , \FrameAddressRegister[14] , \FrameAddressRegister[13] , \FrameAddressRegister[12] , \FrameAddressRegister[11] , \FrameAddressRegister[10] , \FrameAddressRegister[9] , \FrameAddressRegister[8] , \FrameAddressRegister[7] , \FrameAddressRegister[6] , \FrameAddressRegister[5] , \FrameAddressRegister[4] , \FrameAddressRegister[3] , \FrameAddressRegister[2] , \FrameAddressRegister[1] , \FrameAddressRegister[0]  }),
    .FrameStrobe_O({ \FrameSelect[99] , \FrameSelect[98] , \FrameSelect[97] , \FrameSelect[96] , \FrameSelect[95] , \FrameSelect[94] , \FrameSelect[93] , \FrameSelect[92] , \FrameSelect[91] , \FrameSelect[90] , \FrameSelect[89] , \FrameSelect[88] , \FrameSelect[87] , \FrameSelect[86] , \FrameSelect[85] , \FrameSelect[84] , \FrameSelect[83] , \FrameSelect[82] , \FrameSelect[81] , \FrameSelect[80]  })
  );
  Frame_Select_5 Inst_Frame_Select_5 (
    .FrameSelect({ \FrameAddressRegister[31] , \FrameAddressRegister[30] , \FrameAddressRegister[29] , \FrameAddressRegister[28] , \FrameAddressRegister[27]  }),
    .FrameStrobe(LongFrameStrobe),
    .FrameStrobe_I({ \FrameAddressRegister[19] , \FrameAddressRegister[18] , \FrameAddressRegister[17] , \FrameAddressRegister[16] , \FrameAddressRegister[15] , \FrameAddressRegister[14] , \FrameAddressRegister[13] , \FrameAddressRegister[12] , \FrameAddressRegister[11] , \FrameAddressRegister[10] , \FrameAddressRegister[9] , \FrameAddressRegister[8] , \FrameAddressRegister[7] , \FrameAddressRegister[6] , \FrameAddressRegister[5] , \FrameAddressRegister[4] , \FrameAddressRegister[3] , \FrameAddressRegister[2] , \FrameAddressRegister[1] , \FrameAddressRegister[0]  }),
    .FrameStrobe_O({ \FrameSelect[119] , \FrameSelect[118] , \FrameSelect[117] , \FrameSelect[116] , \FrameSelect[115] , \FrameSelect[114] , \FrameSelect[113] , \FrameSelect[112] , \FrameSelect[111] , \FrameSelect[110] , \FrameSelect[109] , \FrameSelect[108] , \FrameSelect[107] , \FrameSelect[106] , \FrameSelect[105] , \FrameSelect[104] , \FrameSelect[103] , \FrameSelect[102] , \FrameSelect[101] , \FrameSelect[100]  })
  );
  Frame_Select_6 Inst_Frame_Select_6 (
    .FrameSelect({ \FrameAddressRegister[31] , \FrameAddressRegister[30] , \FrameAddressRegister[29] , \FrameAddressRegister[28] , \FrameAddressRegister[27]  }),
    .FrameStrobe(LongFrameStrobe),
    .FrameStrobe_I({ \FrameAddressRegister[19] , \FrameAddressRegister[18] , \FrameAddressRegister[17] , \FrameAddressRegister[16] , \FrameAddressRegister[15] , \FrameAddressRegister[14] , \FrameAddressRegister[13] , \FrameAddressRegister[12] , \FrameAddressRegister[11] , \FrameAddressRegister[10] , \FrameAddressRegister[9] , \FrameAddressRegister[8] , \FrameAddressRegister[7] , \FrameAddressRegister[6] , \FrameAddressRegister[5] , \FrameAddressRegister[4] , \FrameAddressRegister[3] , \FrameAddressRegister[2] , \FrameAddressRegister[1] , \FrameAddressRegister[0]  }),
    .FrameStrobe_O({ \FrameSelect[139] , \FrameSelect[138] , \FrameSelect[137] , \FrameSelect[136] , \FrameSelect[135] , \FrameSelect[134] , \FrameSelect[133] , \FrameSelect[132] , \FrameSelect[131] , \FrameSelect[130] , \FrameSelect[129] , \FrameSelect[128] , \FrameSelect[127] , \FrameSelect[126] , \FrameSelect[125] , \FrameSelect[124] , \FrameSelect[123] , \FrameSelect[122] , \FrameSelect[121] , \FrameSelect[120]  })
  );
  Frame_Select_7 Inst_Frame_Select_7 (
    .FrameSelect({ \FrameAddressRegister[31] , \FrameAddressRegister[30] , \FrameAddressRegister[29] , \FrameAddressRegister[28] , \FrameAddressRegister[27]  }),
    .FrameStrobe(LongFrameStrobe),
    .FrameStrobe_I({ \FrameAddressRegister[19] , \FrameAddressRegister[18] , \FrameAddressRegister[17] , \FrameAddressRegister[16] , \FrameAddressRegister[15] , \FrameAddressRegister[14] , \FrameAddressRegister[13] , \FrameAddressRegister[12] , \FrameAddressRegister[11] , \FrameAddressRegister[10] , \FrameAddressRegister[9] , \FrameAddressRegister[8] , \FrameAddressRegister[7] , \FrameAddressRegister[6] , \FrameAddressRegister[5] , \FrameAddressRegister[4] , \FrameAddressRegister[3] , \FrameAddressRegister[2] , \FrameAddressRegister[1] , \FrameAddressRegister[0]  }),
    .FrameStrobe_O({ \FrameSelect[159] , \FrameSelect[158] , \FrameSelect[157] , \FrameSelect[156] , \FrameSelect[155] , \FrameSelect[154] , \FrameSelect[153] , \FrameSelect[152] , \FrameSelect[151] , \FrameSelect[150] , \FrameSelect[149] , \FrameSelect[148] , \FrameSelect[147] , \FrameSelect[146] , \FrameSelect[145] , \FrameSelect[144] , \FrameSelect[143] , \FrameSelect[142] , \FrameSelect[141] , \FrameSelect[140]  })
  );
  Frame_Select_8 Inst_Frame_Select_8 (
    .FrameSelect({ \FrameAddressRegister[31] , \FrameAddressRegister[30] , \FrameAddressRegister[29] , \FrameAddressRegister[28] , \FrameAddressRegister[27]  }),
    .FrameStrobe(LongFrameStrobe),
    .FrameStrobe_I({ \FrameAddressRegister[19] , \FrameAddressRegister[18] , \FrameAddressRegister[17] , \FrameAddressRegister[16] , \FrameAddressRegister[15] , \FrameAddressRegister[14] , \FrameAddressRegister[13] , \FrameAddressRegister[12] , \FrameAddressRegister[11] , \FrameAddressRegister[10] , \FrameAddressRegister[9] , \FrameAddressRegister[8] , \FrameAddressRegister[7] , \FrameAddressRegister[6] , \FrameAddressRegister[5] , \FrameAddressRegister[4] , \FrameAddressRegister[3] , \FrameAddressRegister[2] , \FrameAddressRegister[1] , \FrameAddressRegister[0]  }),
    .FrameStrobe_O({ \FrameSelect[179] , \FrameSelect[178] , \FrameSelect[177] , \FrameSelect[176] , \FrameSelect[175] , \FrameSelect[174] , \FrameSelect[173] , \FrameSelect[172] , \FrameSelect[171] , \FrameSelect[170] , \FrameSelect[169] , \FrameSelect[168] , \FrameSelect[167] , \FrameSelect[166] , \FrameSelect[165] , \FrameSelect[164] , \FrameSelect[163] , \FrameSelect[162] , \FrameSelect[161] , \FrameSelect[160]  })
  );
  Frame_Select_9 Inst_Frame_Select_9 (
    .FrameSelect({ \FrameAddressRegister[31] , \FrameAddressRegister[30] , \FrameAddressRegister[29] , \FrameAddressRegister[28] , \FrameAddressRegister[27]  }),
    .FrameStrobe(LongFrameStrobe),
    .FrameStrobe_I({ \FrameAddressRegister[19] , \FrameAddressRegister[18] , \FrameAddressRegister[17] , \FrameAddressRegister[16] , \FrameAddressRegister[15] , \FrameAddressRegister[14] , \FrameAddressRegister[13] , \FrameAddressRegister[12] , \FrameAddressRegister[11] , \FrameAddressRegister[10] , \FrameAddressRegister[9] , \FrameAddressRegister[8] , \FrameAddressRegister[7] , \FrameAddressRegister[6] , \FrameAddressRegister[5] , \FrameAddressRegister[4] , \FrameAddressRegister[3] , \FrameAddressRegister[2] , \FrameAddressRegister[1] , \FrameAddressRegister[0]  }),
    .FrameStrobe_O({ \FrameSelect[199] , \FrameSelect[198] , \FrameSelect[197] , \FrameSelect[196] , \FrameSelect[195] , \FrameSelect[194] , \FrameSelect[193] , \FrameSelect[192] , \FrameSelect[191] , \FrameSelect[190] , \FrameSelect[189] , \FrameSelect[188] , \FrameSelect[187] , \FrameSelect[186] , \FrameSelect[185] , \FrameSelect[184] , \FrameSelect[183] , \FrameSelect[182] , \FrameSelect[181] , \FrameSelect[180]  })
  );
  eFPGA Inst_eFPGA (
    .FrameData({ _074_, _073_, _072_, _036_, _071_, _070_, _035_, _069_, _068_, _067_, _034_, _033_, _066_, _032_, _065_, _064_, _063_, _031_, _062_, _030_, _061_, _029_, _028_, _060_, _059_, _027_, _026_, _025_, _024_, _058_, _057_, _056_, \FrameData[479] , \FrameData[478] , \FrameData[477] , \FrameData[476] , \FrameData[475] , \FrameData[474] , \FrameData[473] , \FrameData[472] , \FrameData[471] , \FrameData[470] , \FrameData[469] , \FrameData[468] , \FrameData[467] , \FrameData[466] , \FrameData[465] , \FrameData[464] , \FrameData[463] , \FrameData[462] , \FrameData[461] , \FrameData[460] , \FrameData[459] , \FrameData[458] , \FrameData[457] , \FrameData[456] , \FrameData[455] , \FrameData[454] , \FrameData[453] , \FrameData[452] , \FrameData[451] , \FrameData[450] , \FrameData[449] , \FrameData[448] , \FrameData[447] , \FrameData[446] , \FrameData[445] , \FrameData[444] , \FrameData[443] , \FrameData[442] , \FrameData[441] , \FrameData[440] , \FrameData[439] , \FrameData[438] , \FrameData[437] , \FrameData[436] , \FrameData[435] , \FrameData[434] , \FrameData[433] , \FrameData[432] , \FrameData[431] , \FrameData[430] , \FrameData[429] , \FrameData[428] , \FrameData[427] , \FrameData[426] , \FrameData[425] , \FrameData[424] , \FrameData[423] , \FrameData[422] , \FrameData[421] , \FrameData[420] , \FrameData[419] , \FrameData[418] , \FrameData[417] , \FrameData[416] , \FrameData[415] , \FrameData[414] , \FrameData[413] , \FrameData[412] , \FrameData[411] , \FrameData[410] , \FrameData[409] , \FrameData[408] , \FrameData[407] , \FrameData[406] , \FrameData[405] , \FrameData[404] , \FrameData[403] , \FrameData[402] , \FrameData[401] , \FrameData[400] , \FrameData[399] , \FrameData[398] , \FrameData[397] , \FrameData[396] , \FrameData[395] , \FrameData[394] , \FrameData[393] , \FrameData[392] , \FrameData[391] , \FrameData[390] , \FrameData[389] , \FrameData[388] , \FrameData[387] , \FrameData[386] , \FrameData[385] , \FrameData[384] , \FrameData[383] , \FrameData[382] , \FrameData[381] , \FrameData[380] , \FrameData[379] , \FrameData[378] , \FrameData[377] , \FrameData[376] , \FrameData[375] , \FrameData[374] , \FrameData[373] , \FrameData[372] , \FrameData[371] , \FrameData[370] , \FrameData[369] , \FrameData[368] , \FrameData[367] , \FrameData[366] , \FrameData[365] , \FrameData[364] , \FrameData[363] , \FrameData[362] , \FrameData[361] , \FrameData[360] , \FrameData[359] , \FrameData[358] , \FrameData[357] , \FrameData[356] , \FrameData[355] , \FrameData[354] , \FrameData[353] , \FrameData[352] , \FrameData[351] , \FrameData[350] , \FrameData[349] , \FrameData[348] , \FrameData[347] , \FrameData[346] , \FrameData[345] , \FrameData[344] , \FrameData[343] , \FrameData[342] , \FrameData[341] , \FrameData[340] , \FrameData[339] , \FrameData[338] , \FrameData[337] , \FrameData[336] , \FrameData[335] , \FrameData[334] , \FrameData[333] , \FrameData[332] , \FrameData[331] , \FrameData[330] , \FrameData[329] , \FrameData[328] , \FrameData[327] , \FrameData[326] , \FrameData[325] , \FrameData[324] , \FrameData[323] , \FrameData[322] , \FrameData[321] , \FrameData[320] , \FrameData[319] , \FrameData[318] , \FrameData[317] , \FrameData[316] , \FrameData[315] , \FrameData[314] , \FrameData[313] , \FrameData[312] , \FrameData[311] , \FrameData[310] , \FrameData[309] , \FrameData[308] , \FrameData[307] , \FrameData[306] , \FrameData[305] , \FrameData[304] , \FrameData[303] , \FrameData[302] , \FrameData[301] , \FrameData[300] , \FrameData[299] , \FrameData[298] , \FrameData[297] , \FrameData[296] , \FrameData[295] , \FrameData[294] , \FrameData[293] , \FrameData[292] , \FrameData[291] , \FrameData[290] , \FrameData[289] , \FrameData[288] , \FrameData[287] , \FrameData[286] , \FrameData[285] , \FrameData[284] , \FrameData[283] , \FrameData[282] , \FrameData[281] , \FrameData[280] , \FrameData[279] , \FrameData[278] , \FrameData[277] , \FrameData[276] , \FrameData[275] , \FrameData[274] , \FrameData[273] , \FrameData[272] , \FrameData[271] , \FrameData[270] , \FrameData[269] , \FrameData[268] , \FrameData[267] , \FrameData[266] , \FrameData[265] , \FrameData[264] , \FrameData[263] , \FrameData[262] , \FrameData[261] , \FrameData[260] , \FrameData[259] , \FrameData[258] , \FrameData[257] , \FrameData[256] , \FrameData[255] , \FrameData[254] , \FrameData[253] , \FrameData[252] , \FrameData[251] , \FrameData[250] , \FrameData[249] , \FrameData[248] , \FrameData[247] , \FrameData[246] , \FrameData[245] , \FrameData[244] , \FrameData[243] , \FrameData[242] , \FrameData[241] , \FrameData[240] , \FrameData[239] , \FrameData[238] , \FrameData[237] , \FrameData[236] , \FrameData[235] , \FrameData[234] , \FrameData[233] , \FrameData[232] , \FrameData[231] , \FrameData[230] , \FrameData[229] , \FrameData[228] , \FrameData[227] , \FrameData[226] , \FrameData[225] , \FrameData[224] , \FrameData[223] , \FrameData[222] , \FrameData[221] , \FrameData[220] , \FrameData[219] , \FrameData[218] , \FrameData[217] , \FrameData[216] , \FrameData[215] , \FrameData[214] , \FrameData[213] , \FrameData[212] , \FrameData[211] , \FrameData[210] , \FrameData[209] , \FrameData[208] , \FrameData[207] , \FrameData[206] , \FrameData[205] , \FrameData[204] , \FrameData[203] , \FrameData[202] , \FrameData[201] , \FrameData[200] , \FrameData[199] , \FrameData[198] , \FrameData[197] , \FrameData[196] , \FrameData[195] , \FrameData[194] , \FrameData[193] , \FrameData[192] , \FrameData[191] , \FrameData[190] , \FrameData[189] , \FrameData[188] , \FrameData[187] , \FrameData[186] , \FrameData[185] , \FrameData[184] , \FrameData[183] , \FrameData[182] , \FrameData[181] , \FrameData[180] , \FrameData[179] , \FrameData[178] , \FrameData[177] , \FrameData[176] , \FrameData[175] , \FrameData[174] , \FrameData[173] , \FrameData[172] , \FrameData[171] , \FrameData[170] , \FrameData[169] , \FrameData[168] , \FrameData[167] , \FrameData[166] , \FrameData[165] , \FrameData[164] , \FrameData[163] , \FrameData[162] , \FrameData[161] , \FrameData[160] , \FrameData[159] , \FrameData[158] , \FrameData[157] , \FrameData[156] , \FrameData[155] , \FrameData[154] , \FrameData[153] , \FrameData[152] , \FrameData[151] , \FrameData[150] , \FrameData[149] , \FrameData[148] , \FrameData[147] , \FrameData[146] , \FrameData[145] , \FrameData[144] , \FrameData[143] , \FrameData[142] , \FrameData[141] , \FrameData[140] , \FrameData[139] , \FrameData[138] , \FrameData[137] , \FrameData[136] , \FrameData[135] , \FrameData[134] , \FrameData[133] , \FrameData[132] , \FrameData[131] , \FrameData[130] , \FrameData[129] , \FrameData[128] , \FrameData[127] , \FrameData[126] , \FrameData[125] , \FrameData[124] , \FrameData[123] , \FrameData[122] , \FrameData[121] , \FrameData[120] , \FrameData[119] , \FrameData[118] , \FrameData[117] , \FrameData[116] , \FrameData[115] , \FrameData[114] , \FrameData[113] , \FrameData[112] , \FrameData[111] , \FrameData[110] , \FrameData[109] , \FrameData[108] , \FrameData[107] , \FrameData[106] , \FrameData[105] , \FrameData[104] , \FrameData[103] , \FrameData[102] , \FrameData[101] , \FrameData[100] , \FrameData[99] , \FrameData[98] , \FrameData[97] , \FrameData[96] , \FrameData[95] , \FrameData[94] , \FrameData[93] , \FrameData[92] , \FrameData[91] , \FrameData[90] , \FrameData[89] , \FrameData[88] , \FrameData[87] , \FrameData[86] , \FrameData[85] , \FrameData[84] , \FrameData[83] , \FrameData[82] , \FrameData[81] , \FrameData[80] , \FrameData[79] , \FrameData[78] , \FrameData[77] , \FrameData[76] , \FrameData[75] , \FrameData[74] , \FrameData[73] , \FrameData[72] , \FrameData[71] , \FrameData[70] , \FrameData[69] , \FrameData[68] , \FrameData[67] , \FrameData[66] , \FrameData[65] , \FrameData[64] , \FrameData[63] , \FrameData[62] , \FrameData[61] , \FrameData[60] , \FrameData[59] , \FrameData[58] , \FrameData[57] , \FrameData[56] , \FrameData[55] , \FrameData[54] , \FrameData[53] , \FrameData[52] , \FrameData[51] , \FrameData[50] , \FrameData[49] , \FrameData[48] , \FrameData[47] , \FrameData[46] , \FrameData[45] , \FrameData[44] , \FrameData[43] , \FrameData[42] , \FrameData[41] , \FrameData[40] , \FrameData[39] , \FrameData[38] , \FrameData[37] , \FrameData[36] , \FrameData[35] , \FrameData[34] , \FrameData[33] , \FrameData[32] , _055_, _054_, _053_, _023_, _052_, _051_, _022_, _050_, _049_, _048_, _021_, _020_, _047_, _019_, _046_, _045_, _044_, _018_, _043_, _017_, _042_, _016_, _015_, _041_, _040_, _014_, _013_, _012_, _011_, _039_, _038_, _037_ }),
    .FrameStrobe({ \FrameSelect[299] , \FrameSelect[298] , \FrameSelect[297] , \FrameSelect[296] , \FrameSelect[295] , \FrameSelect[294] , \FrameSelect[293] , \FrameSelect[292] , \FrameSelect[291] , \FrameSelect[290] , \FrameSelect[289] , \FrameSelect[288] , \FrameSelect[287] , \FrameSelect[286] , \FrameSelect[285] , \FrameSelect[284] , \FrameSelect[283] , \FrameSelect[282] , \FrameSelect[281] , \FrameSelect[280] , \FrameSelect[279] , \FrameSelect[278] , \FrameSelect[277] , \FrameSelect[276] , \FrameSelect[275] , \FrameSelect[274] , \FrameSelect[273] , \FrameSelect[272] , \FrameSelect[271] , \FrameSelect[270] , \FrameSelect[269] , \FrameSelect[268] , \FrameSelect[267] , \FrameSelect[266] , \FrameSelect[265] , \FrameSelect[264] , \FrameSelect[263] , \FrameSelect[262] , \FrameSelect[261] , \FrameSelect[260] , \FrameSelect[259] , \FrameSelect[258] , \FrameSelect[257] , \FrameSelect[256] , \FrameSelect[255] , \FrameSelect[254] , \FrameSelect[253] , \FrameSelect[252] , \FrameSelect[251] , \FrameSelect[250] , \FrameSelect[249] , \FrameSelect[248] , \FrameSelect[247] , \FrameSelect[246] , \FrameSelect[245] , \FrameSelect[244] , \FrameSelect[243] , \FrameSelect[242] , \FrameSelect[241] , \FrameSelect[240] , \FrameSelect[239] , \FrameSelect[238] , \FrameSelect[237] , \FrameSelect[236] , \FrameSelect[235] , \FrameSelect[234] , \FrameSelect[233] , \FrameSelect[232] , \FrameSelect[231] , \FrameSelect[230] , \FrameSelect[229] , \FrameSelect[228] , \FrameSelect[227] , \FrameSelect[226] , \FrameSelect[225] , \FrameSelect[224] , \FrameSelect[223] , \FrameSelect[222] , \FrameSelect[221] , \FrameSelect[220] , \FrameSelect[219] , \FrameSelect[218] , \FrameSelect[217] , \FrameSelect[216] , \FrameSelect[215] , \FrameSelect[214] , \FrameSelect[213] , \FrameSelect[212] , \FrameSelect[211] , \FrameSelect[210] , \FrameSelect[209] , \FrameSelect[208] , \FrameSelect[207] , \FrameSelect[206] , \FrameSelect[205] , \FrameSelect[204] , \FrameSelect[203] , \FrameSelect[202] , \FrameSelect[201] , \FrameSelect[200] , \FrameSelect[199] , \FrameSelect[198] , \FrameSelect[197] , \FrameSelect[196] , \FrameSelect[195] , \FrameSelect[194] , \FrameSelect[193] , \FrameSelect[192] , \FrameSelect[191] , \FrameSelect[190] , \FrameSelect[189] , \FrameSelect[188] , \FrameSelect[187] , \FrameSelect[186] , \FrameSelect[185] , \FrameSelect[184] , \FrameSelect[183] , \FrameSelect[182] , \FrameSelect[181] , \FrameSelect[180] , \FrameSelect[179] , \FrameSelect[178] , \FrameSelect[177] , \FrameSelect[176] , \FrameSelect[175] , \FrameSelect[174] , \FrameSelect[173] , \FrameSelect[172] , \FrameSelect[171] , \FrameSelect[170] , \FrameSelect[169] , \FrameSelect[168] , \FrameSelect[167] , \FrameSelect[166] , \FrameSelect[165] , \FrameSelect[164] , \FrameSelect[163] , \FrameSelect[162] , \FrameSelect[161] , \FrameSelect[160] , \FrameSelect[159] , \FrameSelect[158] , \FrameSelect[157] , \FrameSelect[156] , \FrameSelect[155] , \FrameSelect[154] , \FrameSelect[153] , \FrameSelect[152] , \FrameSelect[151] , \FrameSelect[150] , \FrameSelect[149] , \FrameSelect[148] , \FrameSelect[147] , \FrameSelect[146] , \FrameSelect[145] , \FrameSelect[144] , \FrameSelect[143] , \FrameSelect[142] , \FrameSelect[141] , \FrameSelect[140] , \FrameSelect[139] , \FrameSelect[138] , \FrameSelect[137] , \FrameSelect[136] , \FrameSelect[135] , \FrameSelect[134] , \FrameSelect[133] , \FrameSelect[132] , \FrameSelect[131] , \FrameSelect[130] , \FrameSelect[129] , \FrameSelect[128] , \FrameSelect[127] , \FrameSelect[126] , \FrameSelect[125] , \FrameSelect[124] , \FrameSelect[123] , \FrameSelect[122] , \FrameSelect[121] , \FrameSelect[120] , \FrameSelect[119] , \FrameSelect[118] , \FrameSelect[117] , \FrameSelect[116] , \FrameSelect[115] , \FrameSelect[114] , \FrameSelect[113] , \FrameSelect[112] , \FrameSelect[111] , \FrameSelect[110] , \FrameSelect[109] , \FrameSelect[108] , \FrameSelect[107] , \FrameSelect[106] , \FrameSelect[105] , \FrameSelect[104] , \FrameSelect[103] , \FrameSelect[102] , \FrameSelect[101] , \FrameSelect[100] , \FrameSelect[99] , \FrameSelect[98] , \FrameSelect[97] , \FrameSelect[96] , \FrameSelect[95] , \FrameSelect[94] , \FrameSelect[93] , \FrameSelect[92] , \FrameSelect[91] , \FrameSelect[90] , \FrameSelect[89] , \FrameSelect[88] , \FrameSelect[87] , \FrameSelect[86] , \FrameSelect[85] , \FrameSelect[84] , \FrameSelect[83] , \FrameSelect[82] , \FrameSelect[81] , \FrameSelect[80] , \FrameSelect[79] , \FrameSelect[78] , \FrameSelect[77] , \FrameSelect[76] , \FrameSelect[75] , \FrameSelect[74] , \FrameSelect[73] , \FrameSelect[72] , \FrameSelect[71] , \FrameSelect[70] , \FrameSelect[69] , \FrameSelect[68] , \FrameSelect[67] , \FrameSelect[66] , \FrameSelect[65] , \FrameSelect[64] , \FrameSelect[63] , \FrameSelect[62] , \FrameSelect[61] , \FrameSelect[60] , \FrameSelect[59] , \FrameSelect[58] , \FrameSelect[57] , \FrameSelect[56] , \FrameSelect[55] , \FrameSelect[54] , \FrameSelect[53] , \FrameSelect[52] , \FrameSelect[51] , \FrameSelect[50] , \FrameSelect[49] , \FrameSelect[48] , \FrameSelect[47] , \FrameSelect[46] , \FrameSelect[45] , \FrameSelect[44] , \FrameSelect[43] , \FrameSelect[42] , \FrameSelect[41] , \FrameSelect[40] , \FrameSelect[39] , \FrameSelect[38] , \FrameSelect[37] , \FrameSelect[36] , \FrameSelect[35] , \FrameSelect[34] , \FrameSelect[33] , \FrameSelect[32] , \FrameSelect[31] , \FrameSelect[30] , \FrameSelect[29] , \FrameSelect[28] , \FrameSelect[27] , \FrameSelect[26] , \FrameSelect[25] , \FrameSelect[24] , \FrameSelect[23] , \FrameSelect[22] , \FrameSelect[21] , \FrameSelect[20] , \FrameSelect[19] , \FrameSelect[18] , \FrameSelect[17] , \FrameSelect[16] , \FrameSelect[15] , \FrameSelect[14] , \FrameSelect[13] , \FrameSelect[12] , \FrameSelect[11] , \FrameSelect[10] , \FrameSelect[9] , \FrameSelect[8] , \FrameSelect[7] , \FrameSelect[6] , \FrameSelect[5] , \FrameSelect[4] , \FrameSelect[3] , \FrameSelect[2] , \FrameSelect[1] , \FrameSelect[0]  }),
    .Tile_X0Y10_A_I_top(io_out[26]),
    .Tile_X0Y10_A_O_top(io_in[26]),
    .Tile_X0Y10_A_T_top(io_oeb[26]),
    .Tile_X0Y10_A_config_C_bit0(\A_config_C[19] ),
    .Tile_X0Y10_A_config_C_bit1(\A_config_C[18] ),
    .Tile_X0Y10_A_config_C_bit2(\A_config_C[17] ),
    .Tile_X0Y10_A_config_C_bit3(\A_config_C[16] ),
    .Tile_X0Y10_B_I_top(io_out[25]),
    .Tile_X0Y10_B_O_top(io_in[25]),
    .Tile_X0Y10_B_T_top(io_oeb[25]),
    .Tile_X0Y10_B_config_C_bit0(\B_config_C[19] ),
    .Tile_X0Y10_B_config_C_bit1(\B_config_C[18] ),
    .Tile_X0Y10_B_config_C_bit2(\B_config_C[17] ),
    .Tile_X0Y10_B_config_C_bit3(\B_config_C[16] ),
    .Tile_X0Y11_A_I_top(io_out[24]),
    .Tile_X0Y11_A_O_top(io_in[24]),
    .Tile_X0Y11_A_T_top(io_oeb[24]),
    .Tile_X0Y11_A_config_C_bit0(\A_config_C[15] ),
    .Tile_X0Y11_A_config_C_bit1(\A_config_C[14] ),
    .Tile_X0Y11_A_config_C_bit2(\A_config_C[13] ),
    .Tile_X0Y11_A_config_C_bit3(\A_config_C[12] ),
    .Tile_X0Y11_B_I_top(io_out[23]),
    .Tile_X0Y11_B_O_top(io_in[23]),
    .Tile_X0Y11_B_T_top(io_oeb[23]),
    .Tile_X0Y11_B_config_C_bit0(\B_config_C[15] ),
    .Tile_X0Y11_B_config_C_bit1(\B_config_C[14] ),
    .Tile_X0Y11_B_config_C_bit2(\B_config_C[13] ),
    .Tile_X0Y11_B_config_C_bit3(\B_config_C[12] ),
    .Tile_X0Y12_A_I_top(io_out[22]),
    .Tile_X0Y12_A_O_top(io_in[22]),
    .Tile_X0Y12_A_T_top(io_oeb[22]),
    .Tile_X0Y12_A_config_C_bit0(\A_config_C[11] ),
    .Tile_X0Y12_A_config_C_bit1(\A_config_C[10] ),
    .Tile_X0Y12_A_config_C_bit2(\A_config_C[9] ),
    .Tile_X0Y12_A_config_C_bit3(\A_config_C[8] ),
    .Tile_X0Y12_B_I_top(io_out[21]),
    .Tile_X0Y12_B_O_top(io_in[21]),
    .Tile_X0Y12_B_T_top(io_oeb[21]),
    .Tile_X0Y12_B_config_C_bit0(\B_config_C[11] ),
    .Tile_X0Y12_B_config_C_bit1(\B_config_C[10] ),
    .Tile_X0Y12_B_config_C_bit2(\B_config_C[9] ),
    .Tile_X0Y12_B_config_C_bit3(\B_config_C[8] ),
    .Tile_X0Y13_A_I_top(io_out[20]),
    .Tile_X0Y13_A_O_top(io_in[20]),
    .Tile_X0Y13_A_T_top(io_oeb[20]),
    .Tile_X0Y13_A_config_C_bit0(\A_config_C[7] ),
    .Tile_X0Y13_A_config_C_bit1(\A_config_C[6] ),
    .Tile_X0Y13_A_config_C_bit2(\A_config_C[5] ),
    .Tile_X0Y13_A_config_C_bit3(\A_config_C[4] ),
    .Tile_X0Y13_B_I_top(io_out[19]),
    .Tile_X0Y13_B_O_top(io_in[19]),
    .Tile_X0Y13_B_T_top(io_oeb[19]),
    .Tile_X0Y13_B_config_C_bit0(\B_config_C[7] ),
    .Tile_X0Y13_B_config_C_bit1(\B_config_C[6] ),
    .Tile_X0Y13_B_config_C_bit2(\B_config_C[5] ),
    .Tile_X0Y13_B_config_C_bit3(\B_config_C[4] ),
    .Tile_X0Y14_A_I_top(io_out[18]),
    .Tile_X0Y14_A_O_top(io_in[18]),
    .Tile_X0Y14_A_T_top(io_oeb[18]),
    .Tile_X0Y14_A_config_C_bit0(\A_config_C[3] ),
    .Tile_X0Y14_A_config_C_bit1(\A_config_C[2] ),
    .Tile_X0Y14_A_config_C_bit2(\A_config_C[1] ),
    .Tile_X0Y14_A_config_C_bit3(\A_config_C[0] ),
    .Tile_X0Y14_B_I_top(io_out[17]),
    .Tile_X0Y14_B_O_top(io_in[17]),
    .Tile_X0Y14_B_T_top(io_oeb[17]),
    .Tile_X0Y14_B_config_C_bit0(\B_config_C[3] ),
    .Tile_X0Y14_B_config_C_bit1(\B_config_C[2] ),
    .Tile_X0Y14_B_config_C_bit2(\B_config_C[1] ),
    .Tile_X0Y14_B_config_C_bit3(\B_config_C[0] ),
    .Tile_X11Y1_OPA_I0(\E_OPA[35] ),
    .Tile_X11Y1_OPA_I1(\E_OPA[34] ),
    .Tile_X11Y1_OPA_I2(\E_OPA[33] ),
    .Tile_X11Y1_OPA_I3(\E_OPA[32] ),
    .Tile_X11Y1_OPB_I0(\E_OPB[35] ),
    .Tile_X11Y1_OPB_I1(\E_OPB[34] ),
    .Tile_X11Y1_OPB_I2(\E_OPB[33] ),
    .Tile_X11Y1_OPB_I3(\E_OPB[32] ),
    .Tile_X11Y1_RES0_O0(\E_RES0[35] ),
    .Tile_X11Y1_RES0_O1(\E_RES0[34] ),
    .Tile_X11Y1_RES0_O2(\E_RES0[33] ),
    .Tile_X11Y1_RES0_O3(\E_RES0[32] ),
    .Tile_X11Y1_RES1_O0(\E_RES1[35] ),
    .Tile_X11Y1_RES1_O1(\E_RES1[34] ),
    .Tile_X11Y1_RES1_O2(\E_RES1[33] ),
    .Tile_X11Y1_RES1_O3(\E_RES1[32] ),
    .Tile_X11Y1_RES2_O0(\E_RES2[35] ),
    .Tile_X11Y1_RES2_O1(\E_RES2[34] ),
    .Tile_X11Y1_RES2_O2(\E_RES2[33] ),
    .Tile_X11Y1_RES2_O3(\E_RES2[32] ),
    .Tile_X11Y2_OPA_I0(\E_OPA[31] ),
    .Tile_X11Y2_OPA_I1(\E_OPA[30] ),
    .Tile_X11Y2_OPA_I2(\E_OPA[29] ),
    .Tile_X11Y2_OPA_I3(\E_OPA[28] ),
    .Tile_X11Y2_OPB_I0(\E_OPB[31] ),
    .Tile_X11Y2_OPB_I1(\E_OPB[30] ),
    .Tile_X11Y2_OPB_I2(\E_OPB[29] ),
    .Tile_X11Y2_OPB_I3(\E_OPB[28] ),
    .Tile_X11Y2_RES0_O0(\E_RES0[31] ),
    .Tile_X11Y2_RES0_O1(\E_RES0[30] ),
    .Tile_X11Y2_RES0_O2(\E_RES0[29] ),
    .Tile_X11Y2_RES0_O3(\E_RES0[28] ),
    .Tile_X11Y2_RES1_O0(\E_RES1[31] ),
    .Tile_X11Y2_RES1_O1(\E_RES1[30] ),
    .Tile_X11Y2_RES1_O2(\E_RES1[29] ),
    .Tile_X11Y2_RES1_O3(\E_RES1[28] ),
    .Tile_X11Y2_RES2_O0(\E_RES2[31] ),
    .Tile_X11Y2_RES2_O1(\E_RES2[30] ),
    .Tile_X11Y2_RES2_O2(\E_RES2[29] ),
    .Tile_X11Y2_RES2_O3(\E_RES2[28] ),
    .Tile_X11Y3_OPA_I0(\E_OPA[27] ),
    .Tile_X11Y3_OPA_I1(\E_OPA[26] ),
    .Tile_X11Y3_OPA_I2(\E_OPA[25] ),
    .Tile_X11Y3_OPA_I3(\E_OPA[24] ),
    .Tile_X11Y3_OPB_I0(\E_OPB[27] ),
    .Tile_X11Y3_OPB_I1(\E_OPB[26] ),
    .Tile_X11Y3_OPB_I2(\E_OPB[25] ),
    .Tile_X11Y3_OPB_I3(\E_OPB[24] ),
    .Tile_X11Y3_RES0_O0(\E_RES0[27] ),
    .Tile_X11Y3_RES0_O1(\E_RES0[26] ),
    .Tile_X11Y3_RES0_O2(\E_RES0[25] ),
    .Tile_X11Y3_RES0_O3(\E_RES0[24] ),
    .Tile_X11Y3_RES1_O0(\E_RES1[27] ),
    .Tile_X11Y3_RES1_O1(\E_RES1[26] ),
    .Tile_X11Y3_RES1_O2(\E_RES1[25] ),
    .Tile_X11Y3_RES1_O3(\E_RES1[24] ),
    .Tile_X11Y3_RES2_O0(\E_RES2[27] ),
    .Tile_X11Y3_RES2_O1(\E_RES2[26] ),
    .Tile_X11Y3_RES2_O2(\E_RES2[25] ),
    .Tile_X11Y3_RES2_O3(\E_RES2[24] ),
    .Tile_X11Y4_OPA_I0(\E_OPA[23] ),
    .Tile_X11Y4_OPA_I1(\E_OPA[22] ),
    .Tile_X11Y4_OPA_I2(\E_OPA[21] ),
    .Tile_X11Y4_OPA_I3(\E_OPA[20] ),
    .Tile_X11Y4_OPB_I0(\E_OPB[23] ),
    .Tile_X11Y4_OPB_I1(\E_OPB[22] ),
    .Tile_X11Y4_OPB_I2(\E_OPB[21] ),
    .Tile_X11Y4_OPB_I3(\E_OPB[20] ),
    .Tile_X11Y4_RES0_O0(\E_RES0[23] ),
    .Tile_X11Y4_RES0_O1(\E_RES0[22] ),
    .Tile_X11Y4_RES0_O2(\E_RES0[21] ),
    .Tile_X11Y4_RES0_O3(\E_RES0[20] ),
    .Tile_X11Y4_RES1_O0(\E_RES1[23] ),
    .Tile_X11Y4_RES1_O1(\E_RES1[22] ),
    .Tile_X11Y4_RES1_O2(\E_RES1[21] ),
    .Tile_X11Y4_RES1_O3(\E_RES1[20] ),
    .Tile_X11Y4_RES2_O0(\E_RES2[23] ),
    .Tile_X11Y4_RES2_O1(\E_RES2[22] ),
    .Tile_X11Y4_RES2_O2(\E_RES2[21] ),
    .Tile_X11Y4_RES2_O3(\E_RES2[20] ),
    .Tile_X11Y5_OPA_I0(\E_OPA[19] ),
    .Tile_X11Y5_OPA_I1(\E_OPA[18] ),
    .Tile_X11Y5_OPA_I2(\E_OPA[17] ),
    .Tile_X11Y5_OPA_I3(\E_OPA[16] ),
    .Tile_X11Y5_OPB_I0(\E_OPB[19] ),
    .Tile_X11Y5_OPB_I1(\E_OPB[18] ),
    .Tile_X11Y5_OPB_I2(\E_OPB[17] ),
    .Tile_X11Y5_OPB_I3(\E_OPB[16] ),
    .Tile_X11Y5_RES0_O0(\E_RES0[19] ),
    .Tile_X11Y5_RES0_O1(\E_RES0[18] ),
    .Tile_X11Y5_RES0_O2(\E_RES0[17] ),
    .Tile_X11Y5_RES0_O3(\E_RES0[16] ),
    .Tile_X11Y5_RES1_O0(\E_RES1[19] ),
    .Tile_X11Y5_RES1_O1(\E_RES1[18] ),
    .Tile_X11Y5_RES1_O2(\E_RES1[17] ),
    .Tile_X11Y5_RES1_O3(\E_RES1[16] ),
    .Tile_X11Y5_RES2_O0(\E_RES2[19] ),
    .Tile_X11Y5_RES2_O1(\E_RES2[18] ),
    .Tile_X11Y5_RES2_O2(\E_RES2[17] ),
    .Tile_X11Y5_RES2_O3(\E_RES2[16] ),
    .Tile_X11Y6_OPA_I0(\E_OPA[15] ),
    .Tile_X11Y6_OPA_I1(\E_OPA[14] ),
    .Tile_X11Y6_OPA_I2(\E_OPA[13] ),
    .Tile_X11Y6_OPA_I3(\E_OPA[12] ),
    .Tile_X11Y6_OPB_I0(\E_OPB[15] ),
    .Tile_X11Y6_OPB_I1(\E_OPB[14] ),
    .Tile_X11Y6_OPB_I2(\E_OPB[13] ),
    .Tile_X11Y6_OPB_I3(\E_OPB[12] ),
    .Tile_X11Y6_RES0_O0(\E_RES0[15] ),
    .Tile_X11Y6_RES0_O1(\E_RES0[14] ),
    .Tile_X11Y6_RES0_O2(\E_RES0[13] ),
    .Tile_X11Y6_RES0_O3(\E_RES0[12] ),
    .Tile_X11Y6_RES1_O0(\E_RES1[15] ),
    .Tile_X11Y6_RES1_O1(\E_RES1[14] ),
    .Tile_X11Y6_RES1_O2(\E_RES1[13] ),
    .Tile_X11Y6_RES1_O3(\E_RES1[12] ),
    .Tile_X11Y6_RES2_O0(\E_RES2[15] ),
    .Tile_X11Y6_RES2_O1(\E_RES2[14] ),
    .Tile_X11Y6_RES2_O2(\E_RES2[13] ),
    .Tile_X11Y6_RES2_O3(\E_RES2[12] ),
    .Tile_X11Y7_OPA_I0(\E_OPA[11] ),
    .Tile_X11Y7_OPA_I1(\E_OPA[10] ),
    .Tile_X11Y7_OPA_I2(\E_OPA[9] ),
    .Tile_X11Y7_OPA_I3(\E_OPA[8] ),
    .Tile_X11Y7_OPB_I0(\E_OPB[11] ),
    .Tile_X11Y7_OPB_I1(\E_OPB[10] ),
    .Tile_X11Y7_OPB_I2(\E_OPB[9] ),
    .Tile_X11Y7_OPB_I3(\E_OPB[8] ),
    .Tile_X11Y7_RES0_O0(\E_RES0[11] ),
    .Tile_X11Y7_RES0_O1(\E_RES0[10] ),
    .Tile_X11Y7_RES0_O2(\E_RES0[9] ),
    .Tile_X11Y7_RES0_O3(\E_RES0[8] ),
    .Tile_X11Y7_RES1_O0(\E_RES1[11] ),
    .Tile_X11Y7_RES1_O1(\E_RES1[10] ),
    .Tile_X11Y7_RES1_O2(\E_RES1[9] ),
    .Tile_X11Y7_RES1_O3(\E_RES1[8] ),
    .Tile_X11Y7_RES2_O0(\E_RES2[11] ),
    .Tile_X11Y7_RES2_O1(\E_RES2[10] ),
    .Tile_X11Y7_RES2_O2(\E_RES2[9] ),
    .Tile_X11Y7_RES2_O3(\E_RES2[8] ),
    .Tile_X11Y8_OPA_I0(\E_OPA[7] ),
    .Tile_X11Y8_OPA_I1(\E_OPA[6] ),
    .Tile_X11Y8_OPA_I2(\E_OPA[5] ),
    .Tile_X11Y8_OPA_I3(\E_OPA[4] ),
    .Tile_X11Y8_OPB_I0(\E_OPB[7] ),
    .Tile_X11Y8_OPB_I1(\E_OPB[6] ),
    .Tile_X11Y8_OPB_I2(\E_OPB[5] ),
    .Tile_X11Y8_OPB_I3(\E_OPB[4] ),
    .Tile_X11Y8_RES0_O0(\E_RES0[7] ),
    .Tile_X11Y8_RES0_O1(\E_RES0[6] ),
    .Tile_X11Y8_RES0_O2(\E_RES0[5] ),
    .Tile_X11Y8_RES0_O3(\E_RES0[4] ),
    .Tile_X11Y8_RES1_O0(\E_RES1[7] ),
    .Tile_X11Y8_RES1_O1(\E_RES1[6] ),
    .Tile_X11Y8_RES1_O2(\E_RES1[5] ),
    .Tile_X11Y8_RES1_O3(\E_RES1[4] ),
    .Tile_X11Y8_RES2_O0(\E_RES2[7] ),
    .Tile_X11Y8_RES2_O1(\E_RES2[6] ),
    .Tile_X11Y8_RES2_O2(\E_RES2[5] ),
    .Tile_X11Y8_RES2_O3(\E_RES2[4] ),
    .Tile_X11Y9_OPA_I0(\E_OPA[3] ),
    .Tile_X11Y9_OPA_I1(\E_OPA[2] ),
    .Tile_X11Y9_OPA_I2(\E_OPA[1] ),
    .Tile_X11Y9_OPA_I3(\E_OPA[0] ),
    .Tile_X11Y9_OPB_I0(\E_OPB[3] ),
    .Tile_X11Y9_OPB_I1(\E_OPB[2] ),
    .Tile_X11Y9_OPB_I2(\E_OPB[1] ),
    .Tile_X11Y9_OPB_I3(\E_OPB[0] ),
    .Tile_X11Y9_RES0_O0(\E_RES0[3] ),
    .Tile_X11Y9_RES0_O1(\E_RES0[2] ),
    .Tile_X11Y9_RES0_O2(\E_RES0[1] ),
    .Tile_X11Y9_RES0_O3(\E_RES0[0] ),
    .Tile_X11Y9_RES1_O0(\E_RES1[3] ),
    .Tile_X11Y9_RES1_O1(\E_RES1[2] ),
    .Tile_X11Y9_RES1_O2(\E_RES1[1] ),
    .Tile_X11Y9_RES1_O3(\E_RES1[0] ),
    .Tile_X11Y9_RES2_O0(\E_RES2[3] ),
    .Tile_X11Y9_RES2_O1(\E_RES2[2] ),
    .Tile_X11Y9_RES2_O2(\E_RES2[1] ),
    .Tile_X11Y9_RES2_O3(\E_RES2[0] ),
    .Tile_X14Y10_Config_accessC_bit0(\Config_accessC[19] ),
    .Tile_X14Y10_Config_accessC_bit1(\Config_accessC[18] ),
    .Tile_X14Y10_Config_accessC_bit2(\Config_accessC[17] ),
    .Tile_X14Y10_Config_accessC_bit3(\Config_accessC[16] ),
    .Tile_X14Y10_FAB2RAM_A0_O0(\FAB2RAM_A[39] ),
    .Tile_X14Y10_FAB2RAM_A0_O1(\FAB2RAM_A[38] ),
    .Tile_X14Y10_FAB2RAM_A0_O2(\FAB2RAM_A[37] ),
    .Tile_X14Y10_FAB2RAM_A0_O3(\FAB2RAM_A[36] ),
    .Tile_X14Y10_FAB2RAM_A1_O0(\FAB2RAM_A[35] ),
    .Tile_X14Y10_FAB2RAM_A1_O1(\FAB2RAM_A[34] ),
    .Tile_X14Y10_FAB2RAM_A1_O2(\FAB2RAM_A[33] ),
    .Tile_X14Y10_FAB2RAM_A1_O3(\FAB2RAM_A[32] ),
    .Tile_X14Y10_FAB2RAM_C_O0(\FAB2RAM_C[19] ),
    .Tile_X14Y10_FAB2RAM_C_O1(\FAB2RAM_C[18] ),
    .Tile_X14Y10_FAB2RAM_C_O2(\FAB2RAM_C[17] ),
    .Tile_X14Y10_FAB2RAM_C_O3(\FAB2RAM_C[16] ),
    .Tile_X14Y10_FAB2RAM_D0_O0(\FAB2RAM_D[79] ),
    .Tile_X14Y10_FAB2RAM_D0_O1(\FAB2RAM_D[78] ),
    .Tile_X14Y10_FAB2RAM_D0_O2(\FAB2RAM_D[77] ),
    .Tile_X14Y10_FAB2RAM_D0_O3(\FAB2RAM_D[76] ),
    .Tile_X14Y10_FAB2RAM_D1_O0(\FAB2RAM_D[75] ),
    .Tile_X14Y10_FAB2RAM_D1_O1(\FAB2RAM_D[74] ),
    .Tile_X14Y10_FAB2RAM_D1_O2(\FAB2RAM_D[73] ),
    .Tile_X14Y10_FAB2RAM_D1_O3(\FAB2RAM_D[72] ),
    .Tile_X14Y10_FAB2RAM_D2_O0(\FAB2RAM_D[71] ),
    .Tile_X14Y10_FAB2RAM_D2_O1(\FAB2RAM_D[70] ),
    .Tile_X14Y10_FAB2RAM_D2_O2(\FAB2RAM_D[69] ),
    .Tile_X14Y10_FAB2RAM_D2_O3(\FAB2RAM_D[68] ),
    .Tile_X14Y10_FAB2RAM_D3_O0(\FAB2RAM_D[67] ),
    .Tile_X14Y10_FAB2RAM_D3_O1(\FAB2RAM_D[66] ),
    .Tile_X14Y10_FAB2RAM_D3_O2(\FAB2RAM_D[65] ),
    .Tile_X14Y10_FAB2RAM_D3_O3(\FAB2RAM_D[64] ),
    .Tile_X14Y10_RAM2FAB_D0_I0(_075_),
    .Tile_X14Y10_RAM2FAB_D0_I1(_076_),
    .Tile_X14Y10_RAM2FAB_D0_I2(_077_),
    .Tile_X14Y10_RAM2FAB_D0_I3(_078_),
    .Tile_X14Y10_RAM2FAB_D1_I0(_079_),
    .Tile_X14Y10_RAM2FAB_D1_I1(_080_),
    .Tile_X14Y10_RAM2FAB_D1_I2(_081_),
    .Tile_X14Y10_RAM2FAB_D1_I3(_082_),
    .Tile_X14Y10_RAM2FAB_D2_I0(_083_),
    .Tile_X14Y10_RAM2FAB_D2_I1(_084_),
    .Tile_X14Y10_RAM2FAB_D2_I2(_085_),
    .Tile_X14Y10_RAM2FAB_D2_I3(_086_),
    .Tile_X14Y10_RAM2FAB_D3_I0(_087_),
    .Tile_X14Y10_RAM2FAB_D3_I1(_088_),
    .Tile_X14Y10_RAM2FAB_D3_I2(_089_),
    .Tile_X14Y10_RAM2FAB_D3_I3(_090_),
    .Tile_X14Y11_Config_accessC_bit0(\Config_accessC[15] ),
    .Tile_X14Y11_Config_accessC_bit1(\Config_accessC[14] ),
    .Tile_X14Y11_Config_accessC_bit2(\Config_accessC[13] ),
    .Tile_X14Y11_Config_accessC_bit3(\Config_accessC[12] ),
    .Tile_X14Y11_FAB2RAM_A0_O0(\FAB2RAM_A[31] ),
    .Tile_X14Y11_FAB2RAM_A0_O1(\FAB2RAM_A[30] ),
    .Tile_X14Y11_FAB2RAM_A0_O2(\FAB2RAM_A[29] ),
    .Tile_X14Y11_FAB2RAM_A0_O3(\FAB2RAM_A[28] ),
    .Tile_X14Y11_FAB2RAM_A1_O0(\FAB2RAM_A[27] ),
    .Tile_X14Y11_FAB2RAM_A1_O1(\FAB2RAM_A[26] ),
    .Tile_X14Y11_FAB2RAM_A1_O2(\FAB2RAM_A[25] ),
    .Tile_X14Y11_FAB2RAM_A1_O3(\FAB2RAM_A[24] ),
    .Tile_X14Y11_FAB2RAM_C_O0(\FAB2RAM_C[15] ),
    .Tile_X14Y11_FAB2RAM_C_O1(\FAB2RAM_C[14] ),
    .Tile_X14Y11_FAB2RAM_C_O2(\FAB2RAM_C[13] ),
    .Tile_X14Y11_FAB2RAM_C_O3(\FAB2RAM_C[12] ),
    .Tile_X14Y11_FAB2RAM_D0_O0(\FAB2RAM_D[63] ),
    .Tile_X14Y11_FAB2RAM_D0_O1(\FAB2RAM_D[62] ),
    .Tile_X14Y11_FAB2RAM_D0_O2(\FAB2RAM_D[61] ),
    .Tile_X14Y11_FAB2RAM_D0_O3(\FAB2RAM_D[60] ),
    .Tile_X14Y11_FAB2RAM_D1_O0(\FAB2RAM_D[59] ),
    .Tile_X14Y11_FAB2RAM_D1_O1(\FAB2RAM_D[58] ),
    .Tile_X14Y11_FAB2RAM_D1_O2(\FAB2RAM_D[57] ),
    .Tile_X14Y11_FAB2RAM_D1_O3(\FAB2RAM_D[56] ),
    .Tile_X14Y11_FAB2RAM_D2_O0(\FAB2RAM_D[55] ),
    .Tile_X14Y11_FAB2RAM_D2_O1(\FAB2RAM_D[54] ),
    .Tile_X14Y11_FAB2RAM_D2_O2(\FAB2RAM_D[53] ),
    .Tile_X14Y11_FAB2RAM_D2_O3(\FAB2RAM_D[52] ),
    .Tile_X14Y11_FAB2RAM_D3_O0(\FAB2RAM_D[51] ),
    .Tile_X14Y11_FAB2RAM_D3_O1(\FAB2RAM_D[50] ),
    .Tile_X14Y11_FAB2RAM_D3_O2(\FAB2RAM_D[49] ),
    .Tile_X14Y11_FAB2RAM_D3_O3(\FAB2RAM_D[48] ),
    .Tile_X14Y11_RAM2FAB_D0_I0(_091_),
    .Tile_X14Y11_RAM2FAB_D0_I1(_092_),
    .Tile_X14Y11_RAM2FAB_D0_I2(_093_),
    .Tile_X14Y11_RAM2FAB_D0_I3(_094_),
    .Tile_X14Y11_RAM2FAB_D1_I0(_095_),
    .Tile_X14Y11_RAM2FAB_D1_I1(_096_),
    .Tile_X14Y11_RAM2FAB_D1_I2(_097_),
    .Tile_X14Y11_RAM2FAB_D1_I3(_098_),
    .Tile_X14Y11_RAM2FAB_D2_I0(_099_),
    .Tile_X14Y11_RAM2FAB_D2_I1(_100_),
    .Tile_X14Y11_RAM2FAB_D2_I2(_101_),
    .Tile_X14Y11_RAM2FAB_D2_I3(_102_),
    .Tile_X14Y11_RAM2FAB_D3_I0(_103_),
    .Tile_X14Y11_RAM2FAB_D3_I1(_104_),
    .Tile_X14Y11_RAM2FAB_D3_I2(_105_),
    .Tile_X14Y11_RAM2FAB_D3_I3(_106_),
    .Tile_X14Y12_Config_accessC_bit0(\Config_accessC[11] ),
    .Tile_X14Y12_Config_accessC_bit1(\Config_accessC[10] ),
    .Tile_X14Y12_Config_accessC_bit2(\Config_accessC[9] ),
    .Tile_X14Y12_Config_accessC_bit3(\Config_accessC[8] ),
    .Tile_X14Y12_FAB2RAM_A0_O0(\FAB2RAM_A[23] ),
    .Tile_X14Y12_FAB2RAM_A0_O1(\FAB2RAM_A[22] ),
    .Tile_X14Y12_FAB2RAM_A0_O2(\FAB2RAM_A[21] ),
    .Tile_X14Y12_FAB2RAM_A0_O3(\FAB2RAM_A[20] ),
    .Tile_X14Y12_FAB2RAM_A1_O0(\FAB2RAM_A[19] ),
    .Tile_X14Y12_FAB2RAM_A1_O1(\FAB2RAM_A[18] ),
    .Tile_X14Y12_FAB2RAM_A1_O2(\FAB2RAM_A[17] ),
    .Tile_X14Y12_FAB2RAM_A1_O3(\FAB2RAM_A[16] ),
    .Tile_X14Y12_FAB2RAM_C_O0(\FAB2RAM_C[11] ),
    .Tile_X14Y12_FAB2RAM_C_O1(\FAB2RAM_C[10] ),
    .Tile_X14Y12_FAB2RAM_C_O2(\FAB2RAM_C[9] ),
    .Tile_X14Y12_FAB2RAM_C_O3(\FAB2RAM_C[8] ),
    .Tile_X14Y12_FAB2RAM_D0_O0(\FAB2RAM_D[47] ),
    .Tile_X14Y12_FAB2RAM_D0_O1(\FAB2RAM_D[46] ),
    .Tile_X14Y12_FAB2RAM_D0_O2(\FAB2RAM_D[45] ),
    .Tile_X14Y12_FAB2RAM_D0_O3(\FAB2RAM_D[44] ),
    .Tile_X14Y12_FAB2RAM_D1_O0(\FAB2RAM_D[43] ),
    .Tile_X14Y12_FAB2RAM_D1_O1(\FAB2RAM_D[42] ),
    .Tile_X14Y12_FAB2RAM_D1_O2(\FAB2RAM_D[41] ),
    .Tile_X14Y12_FAB2RAM_D1_O3(\FAB2RAM_D[40] ),
    .Tile_X14Y12_FAB2RAM_D2_O0(\FAB2RAM_D[39] ),
    .Tile_X14Y12_FAB2RAM_D2_O1(\FAB2RAM_D[38] ),
    .Tile_X14Y12_FAB2RAM_D2_O2(\FAB2RAM_D[37] ),
    .Tile_X14Y12_FAB2RAM_D2_O3(\FAB2RAM_D[36] ),
    .Tile_X14Y12_FAB2RAM_D3_O0(\FAB2RAM_D[35] ),
    .Tile_X14Y12_FAB2RAM_D3_O1(\FAB2RAM_D[34] ),
    .Tile_X14Y12_FAB2RAM_D3_O2(\FAB2RAM_D[33] ),
    .Tile_X14Y12_FAB2RAM_D3_O3(\FAB2RAM_D[32] ),
    .Tile_X14Y12_RAM2FAB_D0_I0(_107_),
    .Tile_X14Y12_RAM2FAB_D0_I1(_108_),
    .Tile_X14Y12_RAM2FAB_D0_I2(_109_),
    .Tile_X14Y12_RAM2FAB_D0_I3(_110_),
    .Tile_X14Y12_RAM2FAB_D1_I0(_111_),
    .Tile_X14Y12_RAM2FAB_D1_I1(_112_),
    .Tile_X14Y12_RAM2FAB_D1_I2(_113_),
    .Tile_X14Y12_RAM2FAB_D1_I3(_114_),
    .Tile_X14Y12_RAM2FAB_D2_I0(_115_),
    .Tile_X14Y12_RAM2FAB_D2_I1(_116_),
    .Tile_X14Y12_RAM2FAB_D2_I2(_117_),
    .Tile_X14Y12_RAM2FAB_D2_I3(_118_),
    .Tile_X14Y12_RAM2FAB_D3_I0(_119_),
    .Tile_X14Y12_RAM2FAB_D3_I1(_120_),
    .Tile_X14Y12_RAM2FAB_D3_I2(_121_),
    .Tile_X14Y12_RAM2FAB_D3_I3(_122_),
    .Tile_X14Y13_Config_accessC_bit0(\Config_accessC[7] ),
    .Tile_X14Y13_Config_accessC_bit1(\Config_accessC[6] ),
    .Tile_X14Y13_Config_accessC_bit2(\Config_accessC[5] ),
    .Tile_X14Y13_Config_accessC_bit3(\Config_accessC[4] ),
    .Tile_X14Y13_FAB2RAM_A0_O0(\FAB2RAM_A[15] ),
    .Tile_X14Y13_FAB2RAM_A0_O1(\FAB2RAM_A[14] ),
    .Tile_X14Y13_FAB2RAM_A0_O2(\FAB2RAM_A[13] ),
    .Tile_X14Y13_FAB2RAM_A0_O3(\FAB2RAM_A[12] ),
    .Tile_X14Y13_FAB2RAM_A1_O0(\FAB2RAM_A[11] ),
    .Tile_X14Y13_FAB2RAM_A1_O1(\FAB2RAM_A[10] ),
    .Tile_X14Y13_FAB2RAM_A1_O2(\FAB2RAM_A[9] ),
    .Tile_X14Y13_FAB2RAM_A1_O3(\FAB2RAM_A[8] ),
    .Tile_X14Y13_FAB2RAM_C_O0(\FAB2RAM_C[7] ),
    .Tile_X14Y13_FAB2RAM_C_O1(\FAB2RAM_C[6] ),
    .Tile_X14Y13_FAB2RAM_C_O2(\FAB2RAM_C[5] ),
    .Tile_X14Y13_FAB2RAM_C_O3(\FAB2RAM_C[4] ),
    .Tile_X14Y13_FAB2RAM_D0_O0(\FAB2RAM_D[31] ),
    .Tile_X14Y13_FAB2RAM_D0_O1(\FAB2RAM_D[30] ),
    .Tile_X14Y13_FAB2RAM_D0_O2(\FAB2RAM_D[29] ),
    .Tile_X14Y13_FAB2RAM_D0_O3(\FAB2RAM_D[28] ),
    .Tile_X14Y13_FAB2RAM_D1_O0(\FAB2RAM_D[27] ),
    .Tile_X14Y13_FAB2RAM_D1_O1(\FAB2RAM_D[26] ),
    .Tile_X14Y13_FAB2RAM_D1_O2(\FAB2RAM_D[25] ),
    .Tile_X14Y13_FAB2RAM_D1_O3(\FAB2RAM_D[24] ),
    .Tile_X14Y13_FAB2RAM_D2_O0(\FAB2RAM_D[23] ),
    .Tile_X14Y13_FAB2RAM_D2_O1(\FAB2RAM_D[22] ),
    .Tile_X14Y13_FAB2RAM_D2_O2(\FAB2RAM_D[21] ),
    .Tile_X14Y13_FAB2RAM_D2_O3(\FAB2RAM_D[20] ),
    .Tile_X14Y13_FAB2RAM_D3_O0(\FAB2RAM_D[19] ),
    .Tile_X14Y13_FAB2RAM_D3_O1(\FAB2RAM_D[18] ),
    .Tile_X14Y13_FAB2RAM_D3_O2(\FAB2RAM_D[17] ),
    .Tile_X14Y13_FAB2RAM_D3_O3(\FAB2RAM_D[16] ),
    .Tile_X14Y13_RAM2FAB_D0_I0(_123_),
    .Tile_X14Y13_RAM2FAB_D0_I1(_124_),
    .Tile_X14Y13_RAM2FAB_D0_I2(_125_),
    .Tile_X14Y13_RAM2FAB_D0_I3(_126_),
    .Tile_X14Y13_RAM2FAB_D1_I0(_127_),
    .Tile_X14Y13_RAM2FAB_D1_I1(_128_),
    .Tile_X14Y13_RAM2FAB_D1_I2(_129_),
    .Tile_X14Y13_RAM2FAB_D1_I3(_130_),
    .Tile_X14Y13_RAM2FAB_D2_I0(_131_),
    .Tile_X14Y13_RAM2FAB_D2_I1(_132_),
    .Tile_X14Y13_RAM2FAB_D2_I2(_133_),
    .Tile_X14Y13_RAM2FAB_D2_I3(_134_),
    .Tile_X14Y13_RAM2FAB_D3_I0(_135_),
    .Tile_X14Y13_RAM2FAB_D3_I1(_136_),
    .Tile_X14Y13_RAM2FAB_D3_I2(_137_),
    .Tile_X14Y13_RAM2FAB_D3_I3(_138_),
    .Tile_X14Y14_Config_accessC_bit0(\Config_accessC[3] ),
    .Tile_X14Y14_Config_accessC_bit1(\Config_accessC[2] ),
    .Tile_X14Y14_Config_accessC_bit2(\Config_accessC[1] ),
    .Tile_X14Y14_Config_accessC_bit3(\Config_accessC[0] ),
    .Tile_X14Y14_FAB2RAM_A0_O0(\FAB2RAM_A[7] ),
    .Tile_X14Y14_FAB2RAM_A0_O1(\FAB2RAM_A[6] ),
    .Tile_X14Y14_FAB2RAM_A0_O2(\FAB2RAM_A[5] ),
    .Tile_X14Y14_FAB2RAM_A0_O3(\FAB2RAM_A[4] ),
    .Tile_X14Y14_FAB2RAM_A1_O0(\FAB2RAM_A[3] ),
    .Tile_X14Y14_FAB2RAM_A1_O1(\FAB2RAM_A[2] ),
    .Tile_X14Y14_FAB2RAM_A1_O2(\FAB2RAM_A[1] ),
    .Tile_X14Y14_FAB2RAM_A1_O3(\FAB2RAM_A[0] ),
    .Tile_X14Y14_FAB2RAM_C_O0(\FAB2RAM_C[3] ),
    .Tile_X14Y14_FAB2RAM_C_O1(\FAB2RAM_C[2] ),
    .Tile_X14Y14_FAB2RAM_C_O2(\FAB2RAM_C[1] ),
    .Tile_X14Y14_FAB2RAM_C_O3(\FAB2RAM_C[0] ),
    .Tile_X14Y14_FAB2RAM_D0_O0(\FAB2RAM_D[15] ),
    .Tile_X14Y14_FAB2RAM_D0_O1(\FAB2RAM_D[14] ),
    .Tile_X14Y14_FAB2RAM_D0_O2(\FAB2RAM_D[13] ),
    .Tile_X14Y14_FAB2RAM_D0_O3(\FAB2RAM_D[12] ),
    .Tile_X14Y14_FAB2RAM_D1_O0(\FAB2RAM_D[11] ),
    .Tile_X14Y14_FAB2RAM_D1_O1(\FAB2RAM_D[10] ),
    .Tile_X14Y14_FAB2RAM_D1_O2(\FAB2RAM_D[9] ),
    .Tile_X14Y14_FAB2RAM_D1_O3(\FAB2RAM_D[8] ),
    .Tile_X14Y14_FAB2RAM_D2_O0(\FAB2RAM_D[7] ),
    .Tile_X14Y14_FAB2RAM_D2_O1(\FAB2RAM_D[6] ),
    .Tile_X14Y14_FAB2RAM_D2_O2(\FAB2RAM_D[5] ),
    .Tile_X14Y14_FAB2RAM_D2_O3(\FAB2RAM_D[4] ),
    .Tile_X14Y14_FAB2RAM_D3_O0(\FAB2RAM_D[3] ),
    .Tile_X14Y14_FAB2RAM_D3_O1(\FAB2RAM_D[2] ),
    .Tile_X14Y14_FAB2RAM_D3_O2(\FAB2RAM_D[1] ),
    .Tile_X14Y14_FAB2RAM_D3_O3(\FAB2RAM_D[0] ),
    .Tile_X14Y14_RAM2FAB_D0_I0(_139_),
    .Tile_X14Y14_RAM2FAB_D0_I1(_140_),
    .Tile_X14Y14_RAM2FAB_D0_I2(_141_),
    .Tile_X14Y14_RAM2FAB_D0_I3(_142_),
    .Tile_X14Y14_RAM2FAB_D1_I0(_143_),
    .Tile_X14Y14_RAM2FAB_D1_I1(_144_),
    .Tile_X14Y14_RAM2FAB_D1_I2(_145_),
    .Tile_X14Y14_RAM2FAB_D1_I3(_146_),
    .Tile_X14Y14_RAM2FAB_D2_I0(_147_),
    .Tile_X14Y14_RAM2FAB_D2_I1(_148_),
    .Tile_X14Y14_RAM2FAB_D2_I2(_149_),
    .Tile_X14Y14_RAM2FAB_D2_I3(_150_),
    .Tile_X14Y14_RAM2FAB_D3_I0(_151_),
    .Tile_X14Y14_RAM2FAB_D3_I1(_152_),
    .Tile_X14Y14_RAM2FAB_D3_I2(_153_),
    .Tile_X14Y14_RAM2FAB_D3_I3(_154_),
    .Tile_X3Y1_OPA_I0(\W_OPA[35] ),
    .Tile_X3Y1_OPA_I1(\SelfWriteData[31] ),
    .Tile_X3Y1_OPA_I2(\SelfWriteData[30] ),
    .Tile_X3Y1_OPA_I3(\SelfWriteData[29] ),
    .Tile_X3Y1_OPB_I0(\W_OPB[35] ),
    .Tile_X3Y1_OPB_I1(\W_OPB[34] ),
    .Tile_X3Y1_OPB_I2(\W_OPB[33] ),
    .Tile_X3Y1_OPB_I3(\W_OPB[32] ),
    .Tile_X3Y1_RES0_O0(\W_RES0[35] ),
    .Tile_X3Y1_RES0_O1(\W_RES0[34] ),
    .Tile_X3Y1_RES0_O2(\W_RES0[33] ),
    .Tile_X3Y1_RES0_O3(\W_RES0[32] ),
    .Tile_X3Y1_RES1_O0(\W_RES1[35] ),
    .Tile_X3Y1_RES1_O1(\W_RES1[34] ),
    .Tile_X3Y1_RES1_O2(\W_RES1[33] ),
    .Tile_X3Y1_RES1_O3(\W_RES1[32] ),
    .Tile_X3Y1_RES2_O0(\W_RES2[35] ),
    .Tile_X3Y1_RES2_O1(\W_RES2[34] ),
    .Tile_X3Y1_RES2_O2(\W_RES2[33] ),
    .Tile_X3Y1_RES2_O3(\W_RES2[32] ),
    .Tile_X3Y2_OPA_I0(\SelfWriteData[28] ),
    .Tile_X3Y2_OPA_I1(\SelfWriteData[27] ),
    .Tile_X3Y2_OPA_I2(\SelfWriteData[26] ),
    .Tile_X3Y2_OPA_I3(\SelfWriteData[25] ),
    .Tile_X3Y2_OPB_I0(\W_OPB[31] ),
    .Tile_X3Y2_OPB_I1(\W_OPB[30] ),
    .Tile_X3Y2_OPB_I2(\W_OPB[29] ),
    .Tile_X3Y2_OPB_I3(\W_OPB[28] ),
    .Tile_X3Y2_RES0_O0(\W_RES0[31] ),
    .Tile_X3Y2_RES0_O1(\W_RES0[30] ),
    .Tile_X3Y2_RES0_O2(\W_RES0[29] ),
    .Tile_X3Y2_RES0_O3(\W_RES0[28] ),
    .Tile_X3Y2_RES1_O0(\W_RES1[31] ),
    .Tile_X3Y2_RES1_O1(\W_RES1[30] ),
    .Tile_X3Y2_RES1_O2(\W_RES1[29] ),
    .Tile_X3Y2_RES1_O3(\W_RES1[28] ),
    .Tile_X3Y2_RES2_O0(\W_RES2[31] ),
    .Tile_X3Y2_RES2_O1(\W_RES2[30] ),
    .Tile_X3Y2_RES2_O2(\W_RES2[29] ),
    .Tile_X3Y2_RES2_O3(\W_RES2[28] ),
    .Tile_X3Y3_OPA_I0(\SelfWriteData[24] ),
    .Tile_X3Y3_OPA_I1(\SelfWriteData[23] ),
    .Tile_X3Y3_OPA_I2(\SelfWriteData[22] ),
    .Tile_X3Y3_OPA_I3(\SelfWriteData[21] ),
    .Tile_X3Y3_OPB_I0(\W_OPB[27] ),
    .Tile_X3Y3_OPB_I1(\W_OPB[26] ),
    .Tile_X3Y3_OPB_I2(\W_OPB[25] ),
    .Tile_X3Y3_OPB_I3(\W_OPB[24] ),
    .Tile_X3Y3_RES0_O0(\W_RES0[27] ),
    .Tile_X3Y3_RES0_O1(\W_RES0[26] ),
    .Tile_X3Y3_RES0_O2(\W_RES0[25] ),
    .Tile_X3Y3_RES0_O3(\W_RES0[24] ),
    .Tile_X3Y3_RES1_O0(\W_RES1[27] ),
    .Tile_X3Y3_RES1_O1(\W_RES1[26] ),
    .Tile_X3Y3_RES1_O2(\W_RES1[25] ),
    .Tile_X3Y3_RES1_O3(\W_RES1[24] ),
    .Tile_X3Y3_RES2_O0(\W_RES2[27] ),
    .Tile_X3Y3_RES2_O1(\W_RES2[26] ),
    .Tile_X3Y3_RES2_O2(\W_RES2[25] ),
    .Tile_X3Y3_RES2_O3(\W_RES2[24] ),
    .Tile_X3Y4_OPA_I0(\SelfWriteData[20] ),
    .Tile_X3Y4_OPA_I1(\SelfWriteData[19] ),
    .Tile_X3Y4_OPA_I2(\SelfWriteData[18] ),
    .Tile_X3Y4_OPA_I3(\SelfWriteData[17] ),
    .Tile_X3Y4_OPB_I0(\W_OPB[23] ),
    .Tile_X3Y4_OPB_I1(\W_OPB[22] ),
    .Tile_X3Y4_OPB_I2(\W_OPB[21] ),
    .Tile_X3Y4_OPB_I3(\W_OPB[20] ),
    .Tile_X3Y4_RES0_O0(\W_RES0[23] ),
    .Tile_X3Y4_RES0_O1(\W_RES0[22] ),
    .Tile_X3Y4_RES0_O2(\W_RES0[21] ),
    .Tile_X3Y4_RES0_O3(\W_RES0[20] ),
    .Tile_X3Y4_RES1_O0(\W_RES1[23] ),
    .Tile_X3Y4_RES1_O1(\W_RES1[22] ),
    .Tile_X3Y4_RES1_O2(\W_RES1[21] ),
    .Tile_X3Y4_RES1_O3(\W_RES1[20] ),
    .Tile_X3Y4_RES2_O0(\W_RES2[23] ),
    .Tile_X3Y4_RES2_O1(\W_RES2[22] ),
    .Tile_X3Y4_RES2_O2(\W_RES2[21] ),
    .Tile_X3Y4_RES2_O3(\W_RES2[20] ),
    .Tile_X3Y5_OPA_I0(\SelfWriteData[16] ),
    .Tile_X3Y5_OPA_I1(\SelfWriteData[15] ),
    .Tile_X3Y5_OPA_I2(\SelfWriteData[14] ),
    .Tile_X3Y5_OPA_I3(\SelfWriteData[13] ),
    .Tile_X3Y5_OPB_I0(\W_OPB[19] ),
    .Tile_X3Y5_OPB_I1(\W_OPB[18] ),
    .Tile_X3Y5_OPB_I2(\W_OPB[17] ),
    .Tile_X3Y5_OPB_I3(\W_OPB[16] ),
    .Tile_X3Y5_RES0_O0(\W_RES0[19] ),
    .Tile_X3Y5_RES0_O1(\W_RES0[18] ),
    .Tile_X3Y5_RES0_O2(\W_RES0[17] ),
    .Tile_X3Y5_RES0_O3(\W_RES0[16] ),
    .Tile_X3Y5_RES1_O0(\W_RES1[19] ),
    .Tile_X3Y5_RES1_O1(\W_RES1[18] ),
    .Tile_X3Y5_RES1_O2(\W_RES1[17] ),
    .Tile_X3Y5_RES1_O3(\W_RES1[16] ),
    .Tile_X3Y5_RES2_O0(\W_RES2[19] ),
    .Tile_X3Y5_RES2_O1(\W_RES2[18] ),
    .Tile_X3Y5_RES2_O2(\W_RES2[17] ),
    .Tile_X3Y5_RES2_O3(\W_RES2[16] ),
    .Tile_X3Y6_OPA_I0(\SelfWriteData[12] ),
    .Tile_X3Y6_OPA_I1(\SelfWriteData[11] ),
    .Tile_X3Y6_OPA_I2(\SelfWriteData[10] ),
    .Tile_X3Y6_OPA_I3(\SelfWriteData[9] ),
    .Tile_X3Y6_OPB_I0(\W_OPB[15] ),
    .Tile_X3Y6_OPB_I1(\W_OPB[14] ),
    .Tile_X3Y6_OPB_I2(\W_OPB[13] ),
    .Tile_X3Y6_OPB_I3(\W_OPB[12] ),
    .Tile_X3Y6_RES0_O0(\W_RES0[15] ),
    .Tile_X3Y6_RES0_O1(\W_RES0[14] ),
    .Tile_X3Y6_RES0_O2(\W_RES0[13] ),
    .Tile_X3Y6_RES0_O3(\W_RES0[12] ),
    .Tile_X3Y6_RES1_O0(\W_RES1[15] ),
    .Tile_X3Y6_RES1_O1(\W_RES1[14] ),
    .Tile_X3Y6_RES1_O2(\W_RES1[13] ),
    .Tile_X3Y6_RES1_O3(\W_RES1[12] ),
    .Tile_X3Y6_RES2_O0(\W_RES2[15] ),
    .Tile_X3Y6_RES2_O1(\W_RES2[14] ),
    .Tile_X3Y6_RES2_O2(\W_RES2[13] ),
    .Tile_X3Y6_RES2_O3(\W_RES2[12] ),
    .Tile_X3Y7_OPA_I0(\SelfWriteData[8] ),
    .Tile_X3Y7_OPA_I1(\SelfWriteData[7] ),
    .Tile_X3Y7_OPA_I2(\SelfWriteData[6] ),
    .Tile_X3Y7_OPA_I3(\SelfWriteData[5] ),
    .Tile_X3Y7_OPB_I0(\W_OPB[11] ),
    .Tile_X3Y7_OPB_I1(\W_OPB[10] ),
    .Tile_X3Y7_OPB_I2(\W_OPB[9] ),
    .Tile_X3Y7_OPB_I3(\W_OPB[8] ),
    .Tile_X3Y7_RES0_O0(\W_RES0[11] ),
    .Tile_X3Y7_RES0_O1(\W_RES0[10] ),
    .Tile_X3Y7_RES0_O2(\W_RES0[9] ),
    .Tile_X3Y7_RES0_O3(\W_RES0[8] ),
    .Tile_X3Y7_RES1_O0(\W_RES1[11] ),
    .Tile_X3Y7_RES1_O1(\W_RES1[10] ),
    .Tile_X3Y7_RES1_O2(\W_RES1[9] ),
    .Tile_X3Y7_RES1_O3(\W_RES1[8] ),
    .Tile_X3Y7_RES2_O0(\W_RES2[11] ),
    .Tile_X3Y7_RES2_O1(\W_RES2[10] ),
    .Tile_X3Y7_RES2_O2(\W_RES2[9] ),
    .Tile_X3Y7_RES2_O3(\W_RES2[8] ),
    .Tile_X3Y8_OPA_I0(\SelfWriteData[4] ),
    .Tile_X3Y8_OPA_I1(\SelfWriteData[3] ),
    .Tile_X3Y8_OPA_I2(\SelfWriteData[2] ),
    .Tile_X3Y8_OPA_I3(\SelfWriteData[1] ),
    .Tile_X3Y8_OPB_I0(\W_OPB[7] ),
    .Tile_X3Y8_OPB_I1(\W_OPB[6] ),
    .Tile_X3Y8_OPB_I2(\W_OPB[5] ),
    .Tile_X3Y8_OPB_I3(\W_OPB[4] ),
    .Tile_X3Y8_RES0_O0(\W_RES0[7] ),
    .Tile_X3Y8_RES0_O1(\W_RES0[6] ),
    .Tile_X3Y8_RES0_O2(\W_RES0[5] ),
    .Tile_X3Y8_RES0_O3(\W_RES0[4] ),
    .Tile_X3Y8_RES1_O0(\W_RES1[7] ),
    .Tile_X3Y8_RES1_O1(\W_RES1[6] ),
    .Tile_X3Y8_RES1_O2(\W_RES1[5] ),
    .Tile_X3Y8_RES1_O3(\W_RES1[4] ),
    .Tile_X3Y8_RES2_O0(\W_RES2[7] ),
    .Tile_X3Y8_RES2_O1(\W_RES2[6] ),
    .Tile_X3Y8_RES2_O2(\W_RES2[5] ),
    .Tile_X3Y8_RES2_O3(\W_RES2[4] ),
    .Tile_X3Y9_OPA_I0(\SelfWriteData[0] ),
    .Tile_X3Y9_OPA_I1(\W_OPA[2] ),
    .Tile_X3Y9_OPA_I2(\W_OPA[1] ),
    .Tile_X3Y9_OPA_I3(\W_OPA[0] ),
    .Tile_X3Y9_OPB_I0(\W_OPB[3] ),
    .Tile_X3Y9_OPB_I1(\W_OPB[2] ),
    .Tile_X3Y9_OPB_I2(\W_OPB[1] ),
    .Tile_X3Y9_OPB_I3(\W_OPB[0] ),
    .Tile_X3Y9_RES0_O0(\W_RES0[3] ),
    .Tile_X3Y9_RES0_O1(\W_RES0[2] ),
    .Tile_X3Y9_RES0_O2(\W_RES0[1] ),
    .Tile_X3Y9_RES0_O3(\W_RES0[0] ),
    .Tile_X3Y9_RES1_O0(\W_RES1[3] ),
    .Tile_X3Y9_RES1_O1(\W_RES1[2] ),
    .Tile_X3Y9_RES1_O2(\W_RES1[1] ),
    .Tile_X3Y9_RES1_O3(\W_RES1[0] ),
    .Tile_X3Y9_RES2_O0(\W_RES2[3] ),
    .Tile_X3Y9_RES2_O1(\W_RES2[2] ),
    .Tile_X3Y9_RES2_O2(\W_RES2[1] ),
    .Tile_X3Y9_RES2_O3(\W_RES2[0] ),
    .UserCLK(CLK)
  );
`ifdef NO_SOC
  // faster fabric simulation
  assign SelfWriteData = 32'b0;
  assign SelfWriteStrobe = 1'b0;
  assign E_OPA = 1'b0;
  assign E_OPB = 1'b0;
  assign W_OPA = 1'b0;
  assign W_OPB = 1'b0;
`else
  forte_soc_top forte_soc_top_i (
    .debug_req_1_i(debug_req_1),
    .debug_req_2_i(debug_req_2),
    .eFPGA_delay_1_o({ _007_, _006_, \W_OPB[33] , \W_OPB[32]  }),
    .eFPGA_delay_2_o({ _002_, _001_, \E_OPB[33] , \E_OPB[32]  }),
    .eFPGA_en_1_o(\W_OPA[35] ),
    .eFPGA_en_2_o(\E_OPA[35] ),
    .eFPGA_fpga_done_1_i(\W_RES1[34] ),
    .eFPGA_fpga_done_2_i(\E_RES1[34] ),
    .eFPGA_operand_a_1_o({ \SelfWriteData[31] , \SelfWriteData[30] , \SelfWriteData[29] , \SelfWriteData[28] , \SelfWriteData[27] , \SelfWriteData[26] , \SelfWriteData[25] , \SelfWriteData[24] , \SelfWriteData[23] , \SelfWriteData[22] , \SelfWriteData[21] , \SelfWriteData[20] , \SelfWriteData[19] , \SelfWriteData[18] , \SelfWriteData[17] , \SelfWriteData[16] , \SelfWriteData[15] , \SelfWriteData[14] , \SelfWriteData[13] , \SelfWriteData[12] , \SelfWriteData[11] , \SelfWriteData[10] , \SelfWriteData[9] , \SelfWriteData[8] , \SelfWriteData[7] , \SelfWriteData[6] , \SelfWriteData[5] , \SelfWriteData[4] , \SelfWriteData[3] , \SelfWriteData[2] , \SelfWriteData[1] , \SelfWriteData[0]  }),
    .eFPGA_operand_a_2_o({ \E_OPA[34] , \E_OPA[33] , \E_OPA[32] , \E_OPA[31] , \E_OPA[30] , \E_OPA[29] , \E_OPA[28] , \E_OPA[27] , \E_OPA[26] , \E_OPA[25] , \E_OPA[24] , \E_OPA[23] , \E_OPA[22] , \E_OPA[21] , \E_OPA[20] , \E_OPA[19] , \E_OPA[18] , \E_OPA[17] , \E_OPA[16] , \E_OPA[15] , \E_OPA[14] , \E_OPA[13] , \E_OPA[12] , \E_OPA[11] , \E_OPA[10] , \E_OPA[9] , \E_OPA[8] , \E_OPA[7] , \E_OPA[6] , \E_OPA[5] , \E_OPA[4] , \E_OPA[3]  }),
    .eFPGA_operand_b_1_o({ \W_OPB[31] , \W_OPB[30] , \W_OPB[29] , \W_OPB[28] , \W_OPB[27] , \W_OPB[26] , \W_OPB[25] , \W_OPB[24] , \W_OPB[23] , \W_OPB[22] , \W_OPB[21] , \W_OPB[20] , \W_OPB[19] , \W_OPB[18] , \W_OPB[17] , \W_OPB[16] , \W_OPB[15] , \W_OPB[14] , \W_OPB[13] , \W_OPB[12] , \W_OPB[11] , \W_OPB[10] , \W_OPB[9] , \W_OPB[8] , \W_OPB[7] , \W_OPB[6] , \W_OPB[5] , \W_OPB[4] , \W_OPB[3] , \W_OPB[2] , \W_OPB[1] , \W_OPB[0]  }),
    .eFPGA_operand_b_2_o({ \E_OPB[31] , \E_OPB[30] , \E_OPB[29] , \E_OPB[28] , \E_OPB[27] , \E_OPB[26] , \E_OPB[25] , \E_OPB[24] , \E_OPB[23] , \E_OPB[22] , \E_OPB[21] , \E_OPB[20] , \E_OPB[19] , \E_OPB[18] , \E_OPB[17] , \E_OPB[16] , \E_OPB[15] , \E_OPB[14] , \E_OPB[13] , \E_OPB[12] , \E_OPB[11] , \E_OPB[10] , \E_OPB[9] , \E_OPB[8] , \E_OPB[7] , \E_OPB[6] , \E_OPB[5] , \E_OPB[4] , \E_OPB[3] , \E_OPB[2] , \E_OPB[1] , \E_OPB[0]  }),
    .eFPGA_operator_1_o({ \W_OPB[35] , \W_OPB[34]  }),
    .eFPGA_operator_2_o({ \E_OPB[35] , \E_OPB[34]  }),
    .eFPGA_result_a_1_i({ \W_RES0[31] , \W_RES0[30] , \W_RES0[29] , \W_RES0[28] , \W_RES0[27] , \W_RES0[26] , \W_RES0[25] , \W_RES0[24] , \W_RES0[23] , \W_RES0[22] , \W_RES0[21] , \W_RES0[20] , \W_RES0[19] , \W_RES0[18] , \W_RES0[17] , \W_RES0[16] , \W_RES0[15] , \W_RES0[14] , \W_RES0[13] , \W_RES0[12] , \W_RES0[11] , \W_RES0[10] , \W_RES0[9] , \W_RES0[8] , \W_RES0[7] , \W_RES0[6] , \W_RES0[5] , \W_RES0[4] , \W_RES0[3] , \W_RES0[2] , \W_RES0[1] , \W_RES0[0]  }),
    .eFPGA_result_a_2_i({ \E_RES0[31] , \E_RES0[30] , \E_RES0[29] , \E_RES0[28] , \E_RES0[27] , \E_RES0[26] , \E_RES0[25] , \E_RES0[24] , \E_RES0[23] , \E_RES0[22] , \E_RES0[21] , \E_RES0[20] , \E_RES0[19] , \E_RES0[18] , \E_RES0[17] , \E_RES0[16] , \E_RES0[15] , \E_RES0[14] , \E_RES0[13] , \E_RES0[12] , \E_RES0[11] , \E_RES0[10] , \E_RES0[9] , \E_RES0[8] , \E_RES0[7] , \E_RES0[6] , \E_RES0[5] , \E_RES0[4] , \E_RES0[3] , \E_RES0[2] , \E_RES0[1] , \E_RES0[0]  }),
    .eFPGA_result_b_1_i({ \W_RES1[31] , \W_RES1[30] , \W_RES1[29] , \W_RES1[28] , \W_RES1[27] , \W_RES1[26] , \W_RES1[25] , \W_RES1[24] , \W_RES1[23] , \W_RES1[22] , \W_RES1[21] , \W_RES1[20] , \W_RES1[19] , \W_RES1[18] , \W_RES1[17] , \W_RES1[16] , \W_RES1[15] , \W_RES1[14] , \W_RES1[13] , \W_RES1[12] , \W_RES1[11] , \W_RES1[10] , \W_RES1[9] , \W_RES1[8] , \W_RES1[7] , \W_RES1[6] , \W_RES1[5] , \W_RES1[4] , \W_RES1[3] , \W_RES1[2] , \W_RES1[1] , \W_RES1[0]  }),
    .eFPGA_result_b_2_i({ \E_RES1[31] , \E_RES1[30] , \E_RES1[29] , \E_RES1[28] , \E_RES1[27] , \E_RES1[26] , \E_RES1[25] , \E_RES1[24] , \E_RES1[23] , \E_RES1[22] , \E_RES1[21] , \E_RES1[20] , \E_RES1[19] , \E_RES1[18] , \E_RES1[17] , \E_RES1[16] , \E_RES1[15] , \E_RES1[14] , \E_RES1[13] , \E_RES1[12] , \E_RES1[11] , \E_RES1[10] , \E_RES1[9] , \E_RES1[8] , \E_RES1[7] , \E_RES1[6] , \E_RES1[5] , \E_RES1[4] , \E_RES1[3] , \E_RES1[2] , \E_RES1[1] , \E_RES1[0]  }),
    .eFPGA_result_c_1_i({ \W_RES2[31] , \W_RES2[30] , \W_RES2[29] , \W_RES2[28] , \W_RES2[27] , \W_RES2[26] , \W_RES2[25] , \W_RES2[24] , \W_RES2[23] , \W_RES2[22] , \W_RES2[21] , \W_RES2[20] , \W_RES2[19] , \W_RES2[18] , \W_RES2[17] , \W_RES2[16] , \W_RES2[15] , \W_RES2[14] , \W_RES2[13] , \W_RES2[12] , \W_RES2[11] , \W_RES2[10] , \W_RES2[9] , \W_RES2[8] , \W_RES2[7] , \W_RES2[6] , \W_RES2[5] , \W_RES2[4] , \W_RES2[3] , \W_RES2[2] , \W_RES2[1] , \W_RES2[0]  }),
    .eFPGA_result_c_2_i({ \E_RES2[31] , \E_RES2[30] , \E_RES2[29] , \E_RES2[28] , \E_RES2[27] , \E_RES2[26] , \E_RES2[25] , \E_RES2[24] , \E_RES2[23] , \E_RES2[22] , \E_RES2[21] , \E_RES2[20] , \E_RES2[19] , \E_RES2[18] , \E_RES2[17] , \E_RES2[16] , \E_RES2[15] , \E_RES2[14] , \E_RES2[13] , \E_RES2[12] , \E_RES2[11] , \E_RES2[10] , \E_RES2[9] , \E_RES2[8] , \E_RES2[7] , \E_RES2[6] , \E_RES2[5] , \E_RES2[4] , \E_RES2[3] , \E_RES2[2] , \E_RES2[1] , \E_RES2[0]  }),
    .eFPGA_write_strobe_1_o(SelfWriteStrobe),
    .eFPGA_write_strobe_2_o(io_out[16]),
    .error_uart_to_mem(io_out[16]),
    .fetch_enable_1_i(fetch_enable_1),
    .fetch_enable_2_i(fetch_enable_2),
    .irq_1_i(\W_RES1[33] ),
    .irq_2_i(\E_RES1[33] ),
    .irq_ack_1_o(\W_OPA[0] ),
    .irq_ack_2_o(\E_OPA[0] ),
    .irq_id_1_i({ \W_RES1[32] , \W_RES0[35] , \W_RES0[34] , \W_RES0[33] , \W_RES0[32]  }),
    .irq_id_1_o({ _010_, _009_, _008_, \W_OPA[2] , \W_OPA[1]  }),
    .irq_id_2_i({ \E_RES1[32] , \E_RES0[35] , \E_RES0[34] , \E_RES0[33] , \E_RES0[32]  }),
    .irq_id_2_o({ _005_, _004_, _003_, \E_OPA[2] , \E_OPA[1]  }),
    .rxd_uart(io_in[12]),
    .rxd_uart_to_mem(io_in[14]),
    .txd_uart(io_out[13]),
    .txd_uart_to_mem(io_out[15]),
    .wb_clk_i(CLK),
    .wb_rst_i(wb_rst_i),
    .wbs_ack_o(wbs_ack_o),
    .wbs_adr_i(wbs_adr_i),
    .wbs_cyc_i(wbs_cyc_i),
    .wbs_dat_i(wbs_dat_i),
    .wbs_dat_o(wbs_dat_o),
    .wbs_sel_i(wbs_sel_i),
    .wbs_stb_i(wbs_stb_i),
    .wbs_we_i(wbs_we_i)
  );
`endif
endmodule
