// IMPORTANT NOTE: if using VPR, any instantiated BELs with no outputs MUST be instantiated after IO
// This is because VPR auto-generates names for primitives with no outputs, and we assume OutPass BELs
// are the first BELs to be auto-named in our constraints file.

module template ();
wire Tile_X3Y1_OPA_O0, Tile_X3Y1_OPA_O1, Tile_X3Y1_OPA_O2, Tile_X3Y1_OPA_O3;
(* keep *) InPass4_frame_config Tile_X3Y1_A (.O0(Tile_X3Y1_OPA_O0), .O1(Tile_X3Y1_OPA_O1), .O2(Tile_X3Y1_OPA_O2), .O3(Tile_X3Y1_OPA_O3));

wire Tile_X3Y1_OPB_O0, Tile_X3Y1_OPB_O1, Tile_X3Y1_OPB_O2, Tile_X3Y1_OPB_O3;
(* keep *) InPass4_frame_config Tile_X3Y1_B (.O0(Tile_X3Y1_OPB_O0), .O1(Tile_X3Y1_OPB_O1), .O2(Tile_X3Y1_OPB_O2), .O3(Tile_X3Y1_OPB_O3));

wire Tile_X3Y1_RES0_I0, Tile_X3Y1_RES0_I1, Tile_X3Y1_RES0_I2, Tile_X3Y1_RES0_I3;
(* keep *) OutPass4_frame_config Tile_X3Y1_C (.I0(Tile_X3Y1_RES0_I0), .I1(Tile_X3Y1_RES0_I1), .I2(Tile_X3Y1_RES0_I2), .I3(Tile_X3Y1_RES0_I3));

wire Tile_X3Y1_RES1_I0, Tile_X3Y1_RES1_I1, Tile_X3Y1_RES1_I2, Tile_X3Y1_RES1_I3;
(* keep *) OutPass4_frame_config Tile_X3Y1_D (.I0(Tile_X3Y1_RES1_I0), .I1(Tile_X3Y1_RES1_I1), .I2(Tile_X3Y1_RES1_I2), .I3(Tile_X3Y1_RES1_I3));

wire Tile_X3Y1_RES2_I0, Tile_X3Y1_RES2_I1, Tile_X3Y1_RES2_I2, Tile_X3Y1_RES2_I3;
(* keep *) OutPass4_frame_config Tile_X3Y1_E (.I0(Tile_X3Y1_RES2_I0), .I1(Tile_X3Y1_RES2_I1), .I2(Tile_X3Y1_RES2_I2), .I3(Tile_X3Y1_RES2_I3));

wire Tile_X11Y1_OPA_O0, Tile_X11Y1_OPA_O1, Tile_X11Y1_OPA_O2, Tile_X11Y1_OPA_O3;
(* keep *) InPass4_frame_config Tile_X11Y1_A (.O0(Tile_X11Y1_OPA_O0), .O1(Tile_X11Y1_OPA_O1), .O2(Tile_X11Y1_OPA_O2), .O3(Tile_X11Y1_OPA_O3));

wire Tile_X11Y1_OPB_O0, Tile_X11Y1_OPB_O1, Tile_X11Y1_OPB_O2, Tile_X11Y1_OPB_O3;
(* keep *) InPass4_frame_config Tile_X11Y1_B (.O0(Tile_X11Y1_OPB_O0), .O1(Tile_X11Y1_OPB_O1), .O2(Tile_X11Y1_OPB_O2), .O3(Tile_X11Y1_OPB_O3));

wire Tile_X11Y1_RES0_I0, Tile_X11Y1_RES0_I1, Tile_X11Y1_RES0_I2, Tile_X11Y1_RES0_I3;
(* keep *) OutPass4_frame_config Tile_X11Y1_C (.I0(Tile_X11Y1_RES0_I0), .I1(Tile_X11Y1_RES0_I1), .I2(Tile_X11Y1_RES0_I2), .I3(Tile_X11Y1_RES0_I3));

wire Tile_X11Y1_RES1_I0, Tile_X11Y1_RES1_I1, Tile_X11Y1_RES1_I2, Tile_X11Y1_RES1_I3;
(* keep *) OutPass4_frame_config Tile_X11Y1_D (.I0(Tile_X11Y1_RES1_I0), .I1(Tile_X11Y1_RES1_I1), .I2(Tile_X11Y1_RES1_I2), .I3(Tile_X11Y1_RES1_I3));

wire Tile_X11Y1_RES2_I0, Tile_X11Y1_RES2_I1, Tile_X11Y1_RES2_I2, Tile_X11Y1_RES2_I3;
(* keep *) OutPass4_frame_config Tile_X11Y1_E (.I0(Tile_X11Y1_RES2_I0), .I1(Tile_X11Y1_RES2_I1), .I2(Tile_X11Y1_RES2_I2), .I3(Tile_X11Y1_RES2_I3));

wire Tile_X3Y2_OPA_O0, Tile_X3Y2_OPA_O1, Tile_X3Y2_OPA_O2, Tile_X3Y2_OPA_O3;
(* keep *) InPass4_frame_config Tile_X3Y2_A (.O0(Tile_X3Y2_OPA_O0), .O1(Tile_X3Y2_OPA_O1), .O2(Tile_X3Y2_OPA_O2), .O3(Tile_X3Y2_OPA_O3));

wire Tile_X3Y2_OPB_O0, Tile_X3Y2_OPB_O1, Tile_X3Y2_OPB_O2, Tile_X3Y2_OPB_O3;
(* keep *) InPass4_frame_config Tile_X3Y2_B (.O0(Tile_X3Y2_OPB_O0), .O1(Tile_X3Y2_OPB_O1), .O2(Tile_X3Y2_OPB_O2), .O3(Tile_X3Y2_OPB_O3));

wire Tile_X3Y2_RES0_I0, Tile_X3Y2_RES0_I1, Tile_X3Y2_RES0_I2, Tile_X3Y2_RES0_I3;
(* keep *) OutPass4_frame_config Tile_X3Y2_C (.I0(Tile_X3Y2_RES0_I0), .I1(Tile_X3Y2_RES0_I1), .I2(Tile_X3Y2_RES0_I2), .I3(Tile_X3Y2_RES0_I3));

wire Tile_X3Y2_RES1_I0, Tile_X3Y2_RES1_I1, Tile_X3Y2_RES1_I2, Tile_X3Y2_RES1_I3;
(* keep *) OutPass4_frame_config Tile_X3Y2_D (.I0(Tile_X3Y2_RES1_I0), .I1(Tile_X3Y2_RES1_I1), .I2(Tile_X3Y2_RES1_I2), .I3(Tile_X3Y2_RES1_I3));

wire Tile_X3Y2_RES2_I0, Tile_X3Y2_RES2_I1, Tile_X3Y2_RES2_I2, Tile_X3Y2_RES2_I3;
(* keep *) OutPass4_frame_config Tile_X3Y2_E (.I0(Tile_X3Y2_RES2_I0), .I1(Tile_X3Y2_RES2_I1), .I2(Tile_X3Y2_RES2_I2), .I3(Tile_X3Y2_RES2_I3));

wire Tile_X11Y2_OPA_O0, Tile_X11Y2_OPA_O1, Tile_X11Y2_OPA_O2, Tile_X11Y2_OPA_O3;
(* keep *) InPass4_frame_config Tile_X11Y2_A (.O0(Tile_X11Y2_OPA_O0), .O1(Tile_X11Y2_OPA_O1), .O2(Tile_X11Y2_OPA_O2), .O3(Tile_X11Y2_OPA_O3));

wire Tile_X11Y2_OPB_O0, Tile_X11Y2_OPB_O1, Tile_X11Y2_OPB_O2, Tile_X11Y2_OPB_O3;
(* keep *) InPass4_frame_config Tile_X11Y2_B (.O0(Tile_X11Y2_OPB_O0), .O1(Tile_X11Y2_OPB_O1), .O2(Tile_X11Y2_OPB_O2), .O3(Tile_X11Y2_OPB_O3));

wire Tile_X11Y2_RES0_I0, Tile_X11Y2_RES0_I1, Tile_X11Y2_RES0_I2, Tile_X11Y2_RES0_I3;
(* keep *) OutPass4_frame_config Tile_X11Y2_C (.I0(Tile_X11Y2_RES0_I0), .I1(Tile_X11Y2_RES0_I1), .I2(Tile_X11Y2_RES0_I2), .I3(Tile_X11Y2_RES0_I3));

wire Tile_X11Y2_RES1_I0, Tile_X11Y2_RES1_I1, Tile_X11Y2_RES1_I2, Tile_X11Y2_RES1_I3;
(* keep *) OutPass4_frame_config Tile_X11Y2_D (.I0(Tile_X11Y2_RES1_I0), .I1(Tile_X11Y2_RES1_I1), .I2(Tile_X11Y2_RES1_I2), .I3(Tile_X11Y2_RES1_I3));

wire Tile_X11Y2_RES2_I0, Tile_X11Y2_RES2_I1, Tile_X11Y2_RES2_I2, Tile_X11Y2_RES2_I3;
(* keep *) OutPass4_frame_config Tile_X11Y2_E (.I0(Tile_X11Y2_RES2_I0), .I1(Tile_X11Y2_RES2_I1), .I2(Tile_X11Y2_RES2_I2), .I3(Tile_X11Y2_RES2_I3));

wire Tile_X3Y3_OPA_O0, Tile_X3Y3_OPA_O1, Tile_X3Y3_OPA_O2, Tile_X3Y3_OPA_O3;
(* keep *) InPass4_frame_config Tile_X3Y3_A (.O0(Tile_X3Y3_OPA_O0), .O1(Tile_X3Y3_OPA_O1), .O2(Tile_X3Y3_OPA_O2), .O3(Tile_X3Y3_OPA_O3));

wire Tile_X3Y3_OPB_O0, Tile_X3Y3_OPB_O1, Tile_X3Y3_OPB_O2, Tile_X3Y3_OPB_O3;
(* keep *) InPass4_frame_config Tile_X3Y3_B (.O0(Tile_X3Y3_OPB_O0), .O1(Tile_X3Y3_OPB_O1), .O2(Tile_X3Y3_OPB_O2), .O3(Tile_X3Y3_OPB_O3));

wire Tile_X3Y3_RES0_I0, Tile_X3Y3_RES0_I1, Tile_X3Y3_RES0_I2, Tile_X3Y3_RES0_I3;
(* keep *) OutPass4_frame_config Tile_X3Y3_C (.I0(Tile_X3Y3_RES0_I0), .I1(Tile_X3Y3_RES0_I1), .I2(Tile_X3Y3_RES0_I2), .I3(Tile_X3Y3_RES0_I3));

wire Tile_X3Y3_RES1_I0, Tile_X3Y3_RES1_I1, Tile_X3Y3_RES1_I2, Tile_X3Y3_RES1_I3;
(* keep *) OutPass4_frame_config Tile_X3Y3_D (.I0(Tile_X3Y3_RES1_I0), .I1(Tile_X3Y3_RES1_I1), .I2(Tile_X3Y3_RES1_I2), .I3(Tile_X3Y3_RES1_I3));

wire Tile_X3Y3_RES2_I0, Tile_X3Y3_RES2_I1, Tile_X3Y3_RES2_I2, Tile_X3Y3_RES2_I3;
(* keep *) OutPass4_frame_config Tile_X3Y3_E (.I0(Tile_X3Y3_RES2_I0), .I1(Tile_X3Y3_RES2_I1), .I2(Tile_X3Y3_RES2_I2), .I3(Tile_X3Y3_RES2_I3));

wire Tile_X11Y3_OPA_O0, Tile_X11Y3_OPA_O1, Tile_X11Y3_OPA_O2, Tile_X11Y3_OPA_O3;
(* keep *) InPass4_frame_config Tile_X11Y3_A (.O0(Tile_X11Y3_OPA_O0), .O1(Tile_X11Y3_OPA_O1), .O2(Tile_X11Y3_OPA_O2), .O3(Tile_X11Y3_OPA_O3));

wire Tile_X11Y3_OPB_O0, Tile_X11Y3_OPB_O1, Tile_X11Y3_OPB_O2, Tile_X11Y3_OPB_O3;
(* keep *) InPass4_frame_config Tile_X11Y3_B (.O0(Tile_X11Y3_OPB_O0), .O1(Tile_X11Y3_OPB_O1), .O2(Tile_X11Y3_OPB_O2), .O3(Tile_X11Y3_OPB_O3));

wire Tile_X11Y3_RES0_I0, Tile_X11Y3_RES0_I1, Tile_X11Y3_RES0_I2, Tile_X11Y3_RES0_I3;
(* keep *) OutPass4_frame_config Tile_X11Y3_C (.I0(Tile_X11Y3_RES0_I0), .I1(Tile_X11Y3_RES0_I1), .I2(Tile_X11Y3_RES0_I2), .I3(Tile_X11Y3_RES0_I3));

wire Tile_X11Y3_RES1_I0, Tile_X11Y3_RES1_I1, Tile_X11Y3_RES1_I2, Tile_X11Y3_RES1_I3;
(* keep *) OutPass4_frame_config Tile_X11Y3_D (.I0(Tile_X11Y3_RES1_I0), .I1(Tile_X11Y3_RES1_I1), .I2(Tile_X11Y3_RES1_I2), .I3(Tile_X11Y3_RES1_I3));

wire Tile_X11Y3_RES2_I0, Tile_X11Y3_RES2_I1, Tile_X11Y3_RES2_I2, Tile_X11Y3_RES2_I3;
(* keep *) OutPass4_frame_config Tile_X11Y3_E (.I0(Tile_X11Y3_RES2_I0), .I1(Tile_X11Y3_RES2_I1), .I2(Tile_X11Y3_RES2_I2), .I3(Tile_X11Y3_RES2_I3));

wire Tile_X3Y4_OPA_O0, Tile_X3Y4_OPA_O1, Tile_X3Y4_OPA_O2, Tile_X3Y4_OPA_O3;
(* keep *) InPass4_frame_config Tile_X3Y4_A (.O0(Tile_X3Y4_OPA_O0), .O1(Tile_X3Y4_OPA_O1), .O2(Tile_X3Y4_OPA_O2), .O3(Tile_X3Y4_OPA_O3));

wire Tile_X3Y4_OPB_O0, Tile_X3Y4_OPB_O1, Tile_X3Y4_OPB_O2, Tile_X3Y4_OPB_O3;
(* keep *) InPass4_frame_config Tile_X3Y4_B (.O0(Tile_X3Y4_OPB_O0), .O1(Tile_X3Y4_OPB_O1), .O2(Tile_X3Y4_OPB_O2), .O3(Tile_X3Y4_OPB_O3));

wire Tile_X3Y4_RES0_I0, Tile_X3Y4_RES0_I1, Tile_X3Y4_RES0_I2, Tile_X3Y4_RES0_I3;
(* keep *) OutPass4_frame_config Tile_X3Y4_C (.I0(Tile_X3Y4_RES0_I0), .I1(Tile_X3Y4_RES0_I1), .I2(Tile_X3Y4_RES0_I2), .I3(Tile_X3Y4_RES0_I3));

wire Tile_X3Y4_RES1_I0, Tile_X3Y4_RES1_I1, Tile_X3Y4_RES1_I2, Tile_X3Y4_RES1_I3;
(* keep *) OutPass4_frame_config Tile_X3Y4_D (.I0(Tile_X3Y4_RES1_I0), .I1(Tile_X3Y4_RES1_I1), .I2(Tile_X3Y4_RES1_I2), .I3(Tile_X3Y4_RES1_I3));

wire Tile_X3Y4_RES2_I0, Tile_X3Y4_RES2_I1, Tile_X3Y4_RES2_I2, Tile_X3Y4_RES2_I3;
(* keep *) OutPass4_frame_config Tile_X3Y4_E (.I0(Tile_X3Y4_RES2_I0), .I1(Tile_X3Y4_RES2_I1), .I2(Tile_X3Y4_RES2_I2), .I3(Tile_X3Y4_RES2_I3));

wire Tile_X11Y4_OPA_O0, Tile_X11Y4_OPA_O1, Tile_X11Y4_OPA_O2, Tile_X11Y4_OPA_O3;
(* keep *) InPass4_frame_config Tile_X11Y4_A (.O0(Tile_X11Y4_OPA_O0), .O1(Tile_X11Y4_OPA_O1), .O2(Tile_X11Y4_OPA_O2), .O3(Tile_X11Y4_OPA_O3));

wire Tile_X11Y4_OPB_O0, Tile_X11Y4_OPB_O1, Tile_X11Y4_OPB_O2, Tile_X11Y4_OPB_O3;
(* keep *) InPass4_frame_config Tile_X11Y4_B (.O0(Tile_X11Y4_OPB_O0), .O1(Tile_X11Y4_OPB_O1), .O2(Tile_X11Y4_OPB_O2), .O3(Tile_X11Y4_OPB_O3));

wire Tile_X11Y4_RES0_I0, Tile_X11Y4_RES0_I1, Tile_X11Y4_RES0_I2, Tile_X11Y4_RES0_I3;
(* keep *) OutPass4_frame_config Tile_X11Y4_C (.I0(Tile_X11Y4_RES0_I0), .I1(Tile_X11Y4_RES0_I1), .I2(Tile_X11Y4_RES0_I2), .I3(Tile_X11Y4_RES0_I3));

wire Tile_X11Y4_RES1_I0, Tile_X11Y4_RES1_I1, Tile_X11Y4_RES1_I2, Tile_X11Y4_RES1_I3;
(* keep *) OutPass4_frame_config Tile_X11Y4_D (.I0(Tile_X11Y4_RES1_I0), .I1(Tile_X11Y4_RES1_I1), .I2(Tile_X11Y4_RES1_I2), .I3(Tile_X11Y4_RES1_I3));

wire Tile_X11Y4_RES2_I0, Tile_X11Y4_RES2_I1, Tile_X11Y4_RES2_I2, Tile_X11Y4_RES2_I3;
(* keep *) OutPass4_frame_config Tile_X11Y4_E (.I0(Tile_X11Y4_RES2_I0), .I1(Tile_X11Y4_RES2_I1), .I2(Tile_X11Y4_RES2_I2), .I3(Tile_X11Y4_RES2_I3));

wire Tile_X3Y5_OPA_O0, Tile_X3Y5_OPA_O1, Tile_X3Y5_OPA_O2, Tile_X3Y5_OPA_O3;
(* keep *) InPass4_frame_config Tile_X3Y5_A (.O0(Tile_X3Y5_OPA_O0), .O1(Tile_X3Y5_OPA_O1), .O2(Tile_X3Y5_OPA_O2), .O3(Tile_X3Y5_OPA_O3));

wire Tile_X3Y5_OPB_O0, Tile_X3Y5_OPB_O1, Tile_X3Y5_OPB_O2, Tile_X3Y5_OPB_O3;
(* keep *) InPass4_frame_config Tile_X3Y5_B (.O0(Tile_X3Y5_OPB_O0), .O1(Tile_X3Y5_OPB_O1), .O2(Tile_X3Y5_OPB_O2), .O3(Tile_X3Y5_OPB_O3));

wire Tile_X3Y5_RES0_I0, Tile_X3Y5_RES0_I1, Tile_X3Y5_RES0_I2, Tile_X3Y5_RES0_I3;
(* keep *) OutPass4_frame_config Tile_X3Y5_C (.I0(Tile_X3Y5_RES0_I0), .I1(Tile_X3Y5_RES0_I1), .I2(Tile_X3Y5_RES0_I2), .I3(Tile_X3Y5_RES0_I3));

wire Tile_X3Y5_RES1_I0, Tile_X3Y5_RES1_I1, Tile_X3Y5_RES1_I2, Tile_X3Y5_RES1_I3;
(* keep *) OutPass4_frame_config Tile_X3Y5_D (.I0(Tile_X3Y5_RES1_I0), .I1(Tile_X3Y5_RES1_I1), .I2(Tile_X3Y5_RES1_I2), .I3(Tile_X3Y5_RES1_I3));

wire Tile_X3Y5_RES2_I0, Tile_X3Y5_RES2_I1, Tile_X3Y5_RES2_I2, Tile_X3Y5_RES2_I3;
(* keep *) OutPass4_frame_config Tile_X3Y5_E (.I0(Tile_X3Y5_RES2_I0), .I1(Tile_X3Y5_RES2_I1), .I2(Tile_X3Y5_RES2_I2), .I3(Tile_X3Y5_RES2_I3));

wire Tile_X11Y5_OPA_O0, Tile_X11Y5_OPA_O1, Tile_X11Y5_OPA_O2, Tile_X11Y5_OPA_O3;
(* keep *) InPass4_frame_config Tile_X11Y5_A (.O0(Tile_X11Y5_OPA_O0), .O1(Tile_X11Y5_OPA_O1), .O2(Tile_X11Y5_OPA_O2), .O3(Tile_X11Y5_OPA_O3));

wire Tile_X11Y5_OPB_O0, Tile_X11Y5_OPB_O1, Tile_X11Y5_OPB_O2, Tile_X11Y5_OPB_O3;
(* keep *) InPass4_frame_config Tile_X11Y5_B (.O0(Tile_X11Y5_OPB_O0), .O1(Tile_X11Y5_OPB_O1), .O2(Tile_X11Y5_OPB_O2), .O3(Tile_X11Y5_OPB_O3));

wire Tile_X11Y5_RES0_I0, Tile_X11Y5_RES0_I1, Tile_X11Y5_RES0_I2, Tile_X11Y5_RES0_I3;
(* keep *) OutPass4_frame_config Tile_X11Y5_C (.I0(Tile_X11Y5_RES0_I0), .I1(Tile_X11Y5_RES0_I1), .I2(Tile_X11Y5_RES0_I2), .I3(Tile_X11Y5_RES0_I3));

wire Tile_X11Y5_RES1_I0, Tile_X11Y5_RES1_I1, Tile_X11Y5_RES1_I2, Tile_X11Y5_RES1_I3;
(* keep *) OutPass4_frame_config Tile_X11Y5_D (.I0(Tile_X11Y5_RES1_I0), .I1(Tile_X11Y5_RES1_I1), .I2(Tile_X11Y5_RES1_I2), .I3(Tile_X11Y5_RES1_I3));

wire Tile_X11Y5_RES2_I0, Tile_X11Y5_RES2_I1, Tile_X11Y5_RES2_I2, Tile_X11Y5_RES2_I3;
(* keep *) OutPass4_frame_config Tile_X11Y5_E (.I0(Tile_X11Y5_RES2_I0), .I1(Tile_X11Y5_RES2_I1), .I2(Tile_X11Y5_RES2_I2), .I3(Tile_X11Y5_RES2_I3));

wire Tile_X3Y6_OPA_O0, Tile_X3Y6_OPA_O1, Tile_X3Y6_OPA_O2, Tile_X3Y6_OPA_O3;
(* keep *) InPass4_frame_config Tile_X3Y6_A (.O0(Tile_X3Y6_OPA_O0), .O1(Tile_X3Y6_OPA_O1), .O2(Tile_X3Y6_OPA_O2), .O3(Tile_X3Y6_OPA_O3));

wire Tile_X3Y6_OPB_O0, Tile_X3Y6_OPB_O1, Tile_X3Y6_OPB_O2, Tile_X3Y6_OPB_O3;
(* keep *) InPass4_frame_config Tile_X3Y6_B (.O0(Tile_X3Y6_OPB_O0), .O1(Tile_X3Y6_OPB_O1), .O2(Tile_X3Y6_OPB_O2), .O3(Tile_X3Y6_OPB_O3));

wire Tile_X3Y6_RES0_I0, Tile_X3Y6_RES0_I1, Tile_X3Y6_RES0_I2, Tile_X3Y6_RES0_I3;
(* keep *) OutPass4_frame_config Tile_X3Y6_C (.I0(Tile_X3Y6_RES0_I0), .I1(Tile_X3Y6_RES0_I1), .I2(Tile_X3Y6_RES0_I2), .I3(Tile_X3Y6_RES0_I3));

wire Tile_X3Y6_RES1_I0, Tile_X3Y6_RES1_I1, Tile_X3Y6_RES1_I2, Tile_X3Y6_RES1_I3;
(* keep *) OutPass4_frame_config Tile_X3Y6_D (.I0(Tile_X3Y6_RES1_I0), .I1(Tile_X3Y6_RES1_I1), .I2(Tile_X3Y6_RES1_I2), .I3(Tile_X3Y6_RES1_I3));

wire Tile_X3Y6_RES2_I0, Tile_X3Y6_RES2_I1, Tile_X3Y6_RES2_I2, Tile_X3Y6_RES2_I3;
(* keep *) OutPass4_frame_config Tile_X3Y6_E (.I0(Tile_X3Y6_RES2_I0), .I1(Tile_X3Y6_RES2_I1), .I2(Tile_X3Y6_RES2_I2), .I3(Tile_X3Y6_RES2_I3));

wire Tile_X11Y6_OPA_O0, Tile_X11Y6_OPA_O1, Tile_X11Y6_OPA_O2, Tile_X11Y6_OPA_O3;
(* keep *) InPass4_frame_config Tile_X11Y6_A (.O0(Tile_X11Y6_OPA_O0), .O1(Tile_X11Y6_OPA_O1), .O2(Tile_X11Y6_OPA_O2), .O3(Tile_X11Y6_OPA_O3));

wire Tile_X11Y6_OPB_O0, Tile_X11Y6_OPB_O1, Tile_X11Y6_OPB_O2, Tile_X11Y6_OPB_O3;
(* keep *) InPass4_frame_config Tile_X11Y6_B (.O0(Tile_X11Y6_OPB_O0), .O1(Tile_X11Y6_OPB_O1), .O2(Tile_X11Y6_OPB_O2), .O3(Tile_X11Y6_OPB_O3));

wire Tile_X11Y6_RES0_I0, Tile_X11Y6_RES0_I1, Tile_X11Y6_RES0_I2, Tile_X11Y6_RES0_I3;
(* keep *) OutPass4_frame_config Tile_X11Y6_C (.I0(Tile_X11Y6_RES0_I0), .I1(Tile_X11Y6_RES0_I1), .I2(Tile_X11Y6_RES0_I2), .I3(Tile_X11Y6_RES0_I3));

wire Tile_X11Y6_RES1_I0, Tile_X11Y6_RES1_I1, Tile_X11Y6_RES1_I2, Tile_X11Y6_RES1_I3;
(* keep *) OutPass4_frame_config Tile_X11Y6_D (.I0(Tile_X11Y6_RES1_I0), .I1(Tile_X11Y6_RES1_I1), .I2(Tile_X11Y6_RES1_I2), .I3(Tile_X11Y6_RES1_I3));

wire Tile_X11Y6_RES2_I0, Tile_X11Y6_RES2_I1, Tile_X11Y6_RES2_I2, Tile_X11Y6_RES2_I3;
(* keep *) OutPass4_frame_config Tile_X11Y6_E (.I0(Tile_X11Y6_RES2_I0), .I1(Tile_X11Y6_RES2_I1), .I2(Tile_X11Y6_RES2_I2), .I3(Tile_X11Y6_RES2_I3));

wire Tile_X3Y7_OPA_O0, Tile_X3Y7_OPA_O1, Tile_X3Y7_OPA_O2, Tile_X3Y7_OPA_O3;
(* keep *) InPass4_frame_config Tile_X3Y7_A (.O0(Tile_X3Y7_OPA_O0), .O1(Tile_X3Y7_OPA_O1), .O2(Tile_X3Y7_OPA_O2), .O3(Tile_X3Y7_OPA_O3));

wire Tile_X3Y7_OPB_O0, Tile_X3Y7_OPB_O1, Tile_X3Y7_OPB_O2, Tile_X3Y7_OPB_O3;
(* keep *) InPass4_frame_config Tile_X3Y7_B (.O0(Tile_X3Y7_OPB_O0), .O1(Tile_X3Y7_OPB_O1), .O2(Tile_X3Y7_OPB_O2), .O3(Tile_X3Y7_OPB_O3));

wire Tile_X3Y7_RES0_I0, Tile_X3Y7_RES0_I1, Tile_X3Y7_RES0_I2, Tile_X3Y7_RES0_I3;
(* keep *) OutPass4_frame_config Tile_X3Y7_C (.I0(Tile_X3Y7_RES0_I0), .I1(Tile_X3Y7_RES0_I1), .I2(Tile_X3Y7_RES0_I2), .I3(Tile_X3Y7_RES0_I3));

wire Tile_X3Y7_RES1_I0, Tile_X3Y7_RES1_I1, Tile_X3Y7_RES1_I2, Tile_X3Y7_RES1_I3;
(* keep *) OutPass4_frame_config Tile_X3Y7_D (.I0(Tile_X3Y7_RES1_I0), .I1(Tile_X3Y7_RES1_I1), .I2(Tile_X3Y7_RES1_I2), .I3(Tile_X3Y7_RES1_I3));

wire Tile_X3Y7_RES2_I0, Tile_X3Y7_RES2_I1, Tile_X3Y7_RES2_I2, Tile_X3Y7_RES2_I3;
(* keep *) OutPass4_frame_config Tile_X3Y7_E (.I0(Tile_X3Y7_RES2_I0), .I1(Tile_X3Y7_RES2_I1), .I2(Tile_X3Y7_RES2_I2), .I3(Tile_X3Y7_RES2_I3));

wire Tile_X11Y7_OPA_O0, Tile_X11Y7_OPA_O1, Tile_X11Y7_OPA_O2, Tile_X11Y7_OPA_O3;
(* keep *) InPass4_frame_config Tile_X11Y7_A (.O0(Tile_X11Y7_OPA_O0), .O1(Tile_X11Y7_OPA_O1), .O2(Tile_X11Y7_OPA_O2), .O3(Tile_X11Y7_OPA_O3));

wire Tile_X11Y7_OPB_O0, Tile_X11Y7_OPB_O1, Tile_X11Y7_OPB_O2, Tile_X11Y7_OPB_O3;
(* keep *) InPass4_frame_config Tile_X11Y7_B (.O0(Tile_X11Y7_OPB_O0), .O1(Tile_X11Y7_OPB_O1), .O2(Tile_X11Y7_OPB_O2), .O3(Tile_X11Y7_OPB_O3));

wire Tile_X11Y7_RES0_I0, Tile_X11Y7_RES0_I1, Tile_X11Y7_RES0_I2, Tile_X11Y7_RES0_I3;
(* keep *) OutPass4_frame_config Tile_X11Y7_C (.I0(Tile_X11Y7_RES0_I0), .I1(Tile_X11Y7_RES0_I1), .I2(Tile_X11Y7_RES0_I2), .I3(Tile_X11Y7_RES0_I3));

wire Tile_X11Y7_RES1_I0, Tile_X11Y7_RES1_I1, Tile_X11Y7_RES1_I2, Tile_X11Y7_RES1_I3;
(* keep *) OutPass4_frame_config Tile_X11Y7_D (.I0(Tile_X11Y7_RES1_I0), .I1(Tile_X11Y7_RES1_I1), .I2(Tile_X11Y7_RES1_I2), .I3(Tile_X11Y7_RES1_I3));

wire Tile_X11Y7_RES2_I0, Tile_X11Y7_RES2_I1, Tile_X11Y7_RES2_I2, Tile_X11Y7_RES2_I3;
(* keep *) OutPass4_frame_config Tile_X11Y7_E (.I0(Tile_X11Y7_RES2_I0), .I1(Tile_X11Y7_RES2_I1), .I2(Tile_X11Y7_RES2_I2), .I3(Tile_X11Y7_RES2_I3));

wire Tile_X3Y8_OPA_O0, Tile_X3Y8_OPA_O1, Tile_X3Y8_OPA_O2, Tile_X3Y8_OPA_O3;
(* keep *) InPass4_frame_config Tile_X3Y8_A (.O0(Tile_X3Y8_OPA_O0), .O1(Tile_X3Y8_OPA_O1), .O2(Tile_X3Y8_OPA_O2), .O3(Tile_X3Y8_OPA_O3));

wire Tile_X3Y8_OPB_O0, Tile_X3Y8_OPB_O1, Tile_X3Y8_OPB_O2, Tile_X3Y8_OPB_O3;
(* keep *) InPass4_frame_config Tile_X3Y8_B (.O0(Tile_X3Y8_OPB_O0), .O1(Tile_X3Y8_OPB_O1), .O2(Tile_X3Y8_OPB_O2), .O3(Tile_X3Y8_OPB_O3));

wire Tile_X3Y8_RES0_I0, Tile_X3Y8_RES0_I1, Tile_X3Y8_RES0_I2, Tile_X3Y8_RES0_I3;
(* keep *) OutPass4_frame_config Tile_X3Y8_C (.I0(Tile_X3Y8_RES0_I0), .I1(Tile_X3Y8_RES0_I1), .I2(Tile_X3Y8_RES0_I2), .I3(Tile_X3Y8_RES0_I3));

wire Tile_X3Y8_RES1_I0, Tile_X3Y8_RES1_I1, Tile_X3Y8_RES1_I2, Tile_X3Y8_RES1_I3;
(* keep *) OutPass4_frame_config Tile_X3Y8_D (.I0(Tile_X3Y8_RES1_I0), .I1(Tile_X3Y8_RES1_I1), .I2(Tile_X3Y8_RES1_I2), .I3(Tile_X3Y8_RES1_I3));

wire Tile_X3Y8_RES2_I0, Tile_X3Y8_RES2_I1, Tile_X3Y8_RES2_I2, Tile_X3Y8_RES2_I3;
(* keep *) OutPass4_frame_config Tile_X3Y8_E (.I0(Tile_X3Y8_RES2_I0), .I1(Tile_X3Y8_RES2_I1), .I2(Tile_X3Y8_RES2_I2), .I3(Tile_X3Y8_RES2_I3));

wire Tile_X11Y8_OPA_O0, Tile_X11Y8_OPA_O1, Tile_X11Y8_OPA_O2, Tile_X11Y8_OPA_O3;
(* keep *) InPass4_frame_config Tile_X11Y8_A (.O0(Tile_X11Y8_OPA_O0), .O1(Tile_X11Y8_OPA_O1), .O2(Tile_X11Y8_OPA_O2), .O3(Tile_X11Y8_OPA_O3));

wire Tile_X11Y8_OPB_O0, Tile_X11Y8_OPB_O1, Tile_X11Y8_OPB_O2, Tile_X11Y8_OPB_O3;
(* keep *) InPass4_frame_config Tile_X11Y8_B (.O0(Tile_X11Y8_OPB_O0), .O1(Tile_X11Y8_OPB_O1), .O2(Tile_X11Y8_OPB_O2), .O3(Tile_X11Y8_OPB_O3));

wire Tile_X11Y8_RES0_I0, Tile_X11Y8_RES0_I1, Tile_X11Y8_RES0_I2, Tile_X11Y8_RES0_I3;
(* keep *) OutPass4_frame_config Tile_X11Y8_C (.I0(Tile_X11Y8_RES0_I0), .I1(Tile_X11Y8_RES0_I1), .I2(Tile_X11Y8_RES0_I2), .I3(Tile_X11Y8_RES0_I3));

wire Tile_X11Y8_RES1_I0, Tile_X11Y8_RES1_I1, Tile_X11Y8_RES1_I2, Tile_X11Y8_RES1_I3;
(* keep *) OutPass4_frame_config Tile_X11Y8_D (.I0(Tile_X11Y8_RES1_I0), .I1(Tile_X11Y8_RES1_I1), .I2(Tile_X11Y8_RES1_I2), .I3(Tile_X11Y8_RES1_I3));

wire Tile_X11Y8_RES2_I0, Tile_X11Y8_RES2_I1, Tile_X11Y8_RES2_I2, Tile_X11Y8_RES2_I3;
(* keep *) OutPass4_frame_config Tile_X11Y8_E (.I0(Tile_X11Y8_RES2_I0), .I1(Tile_X11Y8_RES2_I1), .I2(Tile_X11Y8_RES2_I2), .I3(Tile_X11Y8_RES2_I3));

wire Tile_X3Y9_OPA_O0, Tile_X3Y9_OPA_O1, Tile_X3Y9_OPA_O2, Tile_X3Y9_OPA_O3;
(* keep *) InPass4_frame_config Tile_X3Y9_A (.O0(Tile_X3Y9_OPA_O0), .O1(Tile_X3Y9_OPA_O1), .O2(Tile_X3Y9_OPA_O2), .O3(Tile_X3Y9_OPA_O3));

wire Tile_X3Y9_OPB_O0, Tile_X3Y9_OPB_O1, Tile_X3Y9_OPB_O2, Tile_X3Y9_OPB_O3;
(* keep *) InPass4_frame_config Tile_X3Y9_B (.O0(Tile_X3Y9_OPB_O0), .O1(Tile_X3Y9_OPB_O1), .O2(Tile_X3Y9_OPB_O2), .O3(Tile_X3Y9_OPB_O3));

wire Tile_X3Y9_RES0_I0, Tile_X3Y9_RES0_I1, Tile_X3Y9_RES0_I2, Tile_X3Y9_RES0_I3;
(* keep *) OutPass4_frame_config Tile_X3Y9_C (.I0(Tile_X3Y9_RES0_I0), .I1(Tile_X3Y9_RES0_I1), .I2(Tile_X3Y9_RES0_I2), .I3(Tile_X3Y9_RES0_I3));

wire Tile_X3Y9_RES1_I0, Tile_X3Y9_RES1_I1, Tile_X3Y9_RES1_I2, Tile_X3Y9_RES1_I3;
(* keep *) OutPass4_frame_config Tile_X3Y9_D (.I0(Tile_X3Y9_RES1_I0), .I1(Tile_X3Y9_RES1_I1), .I2(Tile_X3Y9_RES1_I2), .I3(Tile_X3Y9_RES1_I3));

wire Tile_X3Y9_RES2_I0, Tile_X3Y9_RES2_I1, Tile_X3Y9_RES2_I2, Tile_X3Y9_RES2_I3;
(* keep *) OutPass4_frame_config Tile_X3Y9_E (.I0(Tile_X3Y9_RES2_I0), .I1(Tile_X3Y9_RES2_I1), .I2(Tile_X3Y9_RES2_I2), .I3(Tile_X3Y9_RES2_I3));

wire Tile_X11Y9_OPA_O0, Tile_X11Y9_OPA_O1, Tile_X11Y9_OPA_O2, Tile_X11Y9_OPA_O3;
(* keep *) InPass4_frame_config Tile_X11Y9_A (.O0(Tile_X11Y9_OPA_O0), .O1(Tile_X11Y9_OPA_O1), .O2(Tile_X11Y9_OPA_O2), .O3(Tile_X11Y9_OPA_O3));

wire Tile_X11Y9_OPB_O0, Tile_X11Y9_OPB_O1, Tile_X11Y9_OPB_O2, Tile_X11Y9_OPB_O3;
(* keep *) InPass4_frame_config Tile_X11Y9_B (.O0(Tile_X11Y9_OPB_O0), .O1(Tile_X11Y9_OPB_O1), .O2(Tile_X11Y9_OPB_O2), .O3(Tile_X11Y9_OPB_O3));

wire Tile_X11Y9_RES0_I0, Tile_X11Y9_RES0_I1, Tile_X11Y9_RES0_I2, Tile_X11Y9_RES0_I3;
(* keep *) OutPass4_frame_config Tile_X11Y9_C (.I0(Tile_X11Y9_RES0_I0), .I1(Tile_X11Y9_RES0_I1), .I2(Tile_X11Y9_RES0_I2), .I3(Tile_X11Y9_RES0_I3));

wire Tile_X11Y9_RES1_I0, Tile_X11Y9_RES1_I1, Tile_X11Y9_RES1_I2, Tile_X11Y9_RES1_I3;
(* keep *) OutPass4_frame_config Tile_X11Y9_D (.I0(Tile_X11Y9_RES1_I0), .I1(Tile_X11Y9_RES1_I1), .I2(Tile_X11Y9_RES1_I2), .I3(Tile_X11Y9_RES1_I3));

wire Tile_X11Y9_RES2_I0, Tile_X11Y9_RES2_I1, Tile_X11Y9_RES2_I2, Tile_X11Y9_RES2_I3;
(* keep *) OutPass4_frame_config Tile_X11Y9_E (.I0(Tile_X11Y9_RES2_I0), .I1(Tile_X11Y9_RES2_I1), .I2(Tile_X11Y9_RES2_I2), .I3(Tile_X11Y9_RES2_I3));

wire Tile_X0Y10_A_I, Tile_X0Y10_A_T, Tile_X0Y10_A_O, Tile_X0Y10_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y10_A (.O(Tile_X0Y10_A_O), .Q(Tile_X0Y10_A_Q), .I(Tile_X0Y10_A_I));

wire Tile_X0Y10_B_I, Tile_X0Y10_B_T, Tile_X0Y10_B_O, Tile_X0Y10_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y10_B (.O(Tile_X0Y10_B_O), .Q(Tile_X0Y10_B_Q), .I(Tile_X0Y10_B_I));

wire Tile_X14Y10_RAM2FAB_D0_O0, Tile_X14Y10_RAM2FAB_D0_O1, Tile_X14Y10_RAM2FAB_D0_O2, Tile_X14Y10_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X14Y10_A (.O0(Tile_X14Y10_RAM2FAB_D0_O0), .O1(Tile_X14Y10_RAM2FAB_D0_O1), .O2(Tile_X14Y10_RAM2FAB_D0_O2), .O3(Tile_X14Y10_RAM2FAB_D0_O3));

wire Tile_X14Y10_RAM2FAB_D1_O0, Tile_X14Y10_RAM2FAB_D1_O1, Tile_X14Y10_RAM2FAB_D1_O2, Tile_X14Y10_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X14Y10_B (.O0(Tile_X14Y10_RAM2FAB_D1_O0), .O1(Tile_X14Y10_RAM2FAB_D1_O1), .O2(Tile_X14Y10_RAM2FAB_D1_O2), .O3(Tile_X14Y10_RAM2FAB_D1_O3));

wire Tile_X14Y10_RAM2FAB_D2_O0, Tile_X14Y10_RAM2FAB_D2_O1, Tile_X14Y10_RAM2FAB_D2_O2, Tile_X14Y10_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X14Y10_C (.O0(Tile_X14Y10_RAM2FAB_D2_O0), .O1(Tile_X14Y10_RAM2FAB_D2_O1), .O2(Tile_X14Y10_RAM2FAB_D2_O2), .O3(Tile_X14Y10_RAM2FAB_D2_O3));

wire Tile_X14Y10_RAM2FAB_D3_O0, Tile_X14Y10_RAM2FAB_D3_O1, Tile_X14Y10_RAM2FAB_D3_O2, Tile_X14Y10_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X14Y10_D (.O0(Tile_X14Y10_RAM2FAB_D3_O0), .O1(Tile_X14Y10_RAM2FAB_D3_O1), .O2(Tile_X14Y10_RAM2FAB_D3_O2), .O3(Tile_X14Y10_RAM2FAB_D3_O3));

wire Tile_X14Y10_FAB2RAM_D0_I0, Tile_X14Y10_FAB2RAM_D0_I1, Tile_X14Y10_FAB2RAM_D0_I2, Tile_X14Y10_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X14Y10_E (.I0(Tile_X14Y10_FAB2RAM_D0_I0), .I1(Tile_X14Y10_FAB2RAM_D0_I1), .I2(Tile_X14Y10_FAB2RAM_D0_I2), .I3(Tile_X14Y10_FAB2RAM_D0_I3));

wire Tile_X14Y10_FAB2RAM_D1_I0, Tile_X14Y10_FAB2RAM_D1_I1, Tile_X14Y10_FAB2RAM_D1_I2, Tile_X14Y10_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X14Y10_F (.I0(Tile_X14Y10_FAB2RAM_D1_I0), .I1(Tile_X14Y10_FAB2RAM_D1_I1), .I2(Tile_X14Y10_FAB2RAM_D1_I2), .I3(Tile_X14Y10_FAB2RAM_D1_I3));

wire Tile_X14Y10_FAB2RAM_D2_I0, Tile_X14Y10_FAB2RAM_D2_I1, Tile_X14Y10_FAB2RAM_D2_I2, Tile_X14Y10_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X14Y10_G (.I0(Tile_X14Y10_FAB2RAM_D2_I0), .I1(Tile_X14Y10_FAB2RAM_D2_I1), .I2(Tile_X14Y10_FAB2RAM_D2_I2), .I3(Tile_X14Y10_FAB2RAM_D2_I3));

wire Tile_X14Y10_FAB2RAM_D3_I0, Tile_X14Y10_FAB2RAM_D3_I1, Tile_X14Y10_FAB2RAM_D3_I2, Tile_X14Y10_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X14Y10_H (.I0(Tile_X14Y10_FAB2RAM_D3_I0), .I1(Tile_X14Y10_FAB2RAM_D3_I1), .I2(Tile_X14Y10_FAB2RAM_D3_I2), .I3(Tile_X14Y10_FAB2RAM_D3_I3));

wire Tile_X14Y10_FAB2RAM_A0_I0, Tile_X14Y10_FAB2RAM_A0_I1, Tile_X14Y10_FAB2RAM_A0_I2, Tile_X14Y10_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X14Y10_I (.I0(Tile_X14Y10_FAB2RAM_A0_I0), .I1(Tile_X14Y10_FAB2RAM_A0_I1), .I2(Tile_X14Y10_FAB2RAM_A0_I2), .I3(Tile_X14Y10_FAB2RAM_A0_I3));

wire Tile_X14Y10_FAB2RAM_A1_I0, Tile_X14Y10_FAB2RAM_A1_I1, Tile_X14Y10_FAB2RAM_A1_I2, Tile_X14Y10_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X14Y10_J (.I0(Tile_X14Y10_FAB2RAM_A1_I0), .I1(Tile_X14Y10_FAB2RAM_A1_I1), .I2(Tile_X14Y10_FAB2RAM_A1_I2), .I3(Tile_X14Y10_FAB2RAM_A1_I3));

wire Tile_X14Y10_FAB2RAM_C_I0, Tile_X14Y10_FAB2RAM_C_I1, Tile_X14Y10_FAB2RAM_C_I2, Tile_X14Y10_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X14Y10_K (.I0(Tile_X14Y10_FAB2RAM_C_I0), .I1(Tile_X14Y10_FAB2RAM_C_I1), .I2(Tile_X14Y10_FAB2RAM_C_I2), .I3(Tile_X14Y10_FAB2RAM_C_I3));

wire Tile_X0Y11_A_I, Tile_X0Y11_A_T, Tile_X0Y11_A_O, Tile_X0Y11_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y11_A (.O(Tile_X0Y11_A_O), .Q(Tile_X0Y11_A_Q), .I(Tile_X0Y11_A_I));

wire Tile_X0Y11_B_I, Tile_X0Y11_B_T, Tile_X0Y11_B_O, Tile_X0Y11_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y11_B (.O(Tile_X0Y11_B_O), .Q(Tile_X0Y11_B_Q), .I(Tile_X0Y11_B_I));

wire Tile_X14Y11_RAM2FAB_D0_O0, Tile_X14Y11_RAM2FAB_D0_O1, Tile_X14Y11_RAM2FAB_D0_O2, Tile_X14Y11_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X14Y11_A (.O0(Tile_X14Y11_RAM2FAB_D0_O0), .O1(Tile_X14Y11_RAM2FAB_D0_O1), .O2(Tile_X14Y11_RAM2FAB_D0_O2), .O3(Tile_X14Y11_RAM2FAB_D0_O3));

wire Tile_X14Y11_RAM2FAB_D1_O0, Tile_X14Y11_RAM2FAB_D1_O1, Tile_X14Y11_RAM2FAB_D1_O2, Tile_X14Y11_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X14Y11_B (.O0(Tile_X14Y11_RAM2FAB_D1_O0), .O1(Tile_X14Y11_RAM2FAB_D1_O1), .O2(Tile_X14Y11_RAM2FAB_D1_O2), .O3(Tile_X14Y11_RAM2FAB_D1_O3));

wire Tile_X14Y11_RAM2FAB_D2_O0, Tile_X14Y11_RAM2FAB_D2_O1, Tile_X14Y11_RAM2FAB_D2_O2, Tile_X14Y11_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X14Y11_C (.O0(Tile_X14Y11_RAM2FAB_D2_O0), .O1(Tile_X14Y11_RAM2FAB_D2_O1), .O2(Tile_X14Y11_RAM2FAB_D2_O2), .O3(Tile_X14Y11_RAM2FAB_D2_O3));

wire Tile_X14Y11_RAM2FAB_D3_O0, Tile_X14Y11_RAM2FAB_D3_O1, Tile_X14Y11_RAM2FAB_D3_O2, Tile_X14Y11_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X14Y11_D (.O0(Tile_X14Y11_RAM2FAB_D3_O0), .O1(Tile_X14Y11_RAM2FAB_D3_O1), .O2(Tile_X14Y11_RAM2FAB_D3_O2), .O3(Tile_X14Y11_RAM2FAB_D3_O3));

wire Tile_X14Y11_FAB2RAM_D0_I0, Tile_X14Y11_FAB2RAM_D0_I1, Tile_X14Y11_FAB2RAM_D0_I2, Tile_X14Y11_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X14Y11_E (.I0(Tile_X14Y11_FAB2RAM_D0_I0), .I1(Tile_X14Y11_FAB2RAM_D0_I1), .I2(Tile_X14Y11_FAB2RAM_D0_I2), .I3(Tile_X14Y11_FAB2RAM_D0_I3));

wire Tile_X14Y11_FAB2RAM_D1_I0, Tile_X14Y11_FAB2RAM_D1_I1, Tile_X14Y11_FAB2RAM_D1_I2, Tile_X14Y11_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X14Y11_F (.I0(Tile_X14Y11_FAB2RAM_D1_I0), .I1(Tile_X14Y11_FAB2RAM_D1_I1), .I2(Tile_X14Y11_FAB2RAM_D1_I2), .I3(Tile_X14Y11_FAB2RAM_D1_I3));

wire Tile_X14Y11_FAB2RAM_D2_I0, Tile_X14Y11_FAB2RAM_D2_I1, Tile_X14Y11_FAB2RAM_D2_I2, Tile_X14Y11_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X14Y11_G (.I0(Tile_X14Y11_FAB2RAM_D2_I0), .I1(Tile_X14Y11_FAB2RAM_D2_I1), .I2(Tile_X14Y11_FAB2RAM_D2_I2), .I3(Tile_X14Y11_FAB2RAM_D2_I3));

wire Tile_X14Y11_FAB2RAM_D3_I0, Tile_X14Y11_FAB2RAM_D3_I1, Tile_X14Y11_FAB2RAM_D3_I2, Tile_X14Y11_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X14Y11_H (.I0(Tile_X14Y11_FAB2RAM_D3_I0), .I1(Tile_X14Y11_FAB2RAM_D3_I1), .I2(Tile_X14Y11_FAB2RAM_D3_I2), .I3(Tile_X14Y11_FAB2RAM_D3_I3));

wire Tile_X14Y11_FAB2RAM_A0_I0, Tile_X14Y11_FAB2RAM_A0_I1, Tile_X14Y11_FAB2RAM_A0_I2, Tile_X14Y11_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X14Y11_I (.I0(Tile_X14Y11_FAB2RAM_A0_I0), .I1(Tile_X14Y11_FAB2RAM_A0_I1), .I2(Tile_X14Y11_FAB2RAM_A0_I2), .I3(Tile_X14Y11_FAB2RAM_A0_I3));

wire Tile_X14Y11_FAB2RAM_A1_I0, Tile_X14Y11_FAB2RAM_A1_I1, Tile_X14Y11_FAB2RAM_A1_I2, Tile_X14Y11_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X14Y11_J (.I0(Tile_X14Y11_FAB2RAM_A1_I0), .I1(Tile_X14Y11_FAB2RAM_A1_I1), .I2(Tile_X14Y11_FAB2RAM_A1_I2), .I3(Tile_X14Y11_FAB2RAM_A1_I3));

wire Tile_X14Y11_FAB2RAM_C_I0, Tile_X14Y11_FAB2RAM_C_I1, Tile_X14Y11_FAB2RAM_C_I2, Tile_X14Y11_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X14Y11_K (.I0(Tile_X14Y11_FAB2RAM_C_I0), .I1(Tile_X14Y11_FAB2RAM_C_I1), .I2(Tile_X14Y11_FAB2RAM_C_I2), .I3(Tile_X14Y11_FAB2RAM_C_I3));

wire Tile_X0Y12_A_I, Tile_X0Y12_A_T, Tile_X0Y12_A_O, Tile_X0Y12_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y12_A (.O(Tile_X0Y12_A_O), .Q(Tile_X0Y12_A_Q), .I(Tile_X0Y12_A_I));

wire Tile_X0Y12_B_I, Tile_X0Y12_B_T, Tile_X0Y12_B_O, Tile_X0Y12_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y12_B (.O(Tile_X0Y12_B_O), .Q(Tile_X0Y12_B_Q), .I(Tile_X0Y12_B_I));

wire Tile_X14Y12_RAM2FAB_D0_O0, Tile_X14Y12_RAM2FAB_D0_O1, Tile_X14Y12_RAM2FAB_D0_O2, Tile_X14Y12_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X14Y12_A (.O0(Tile_X14Y12_RAM2FAB_D0_O0), .O1(Tile_X14Y12_RAM2FAB_D0_O1), .O2(Tile_X14Y12_RAM2FAB_D0_O2), .O3(Tile_X14Y12_RAM2FAB_D0_O3));

wire Tile_X14Y12_RAM2FAB_D1_O0, Tile_X14Y12_RAM2FAB_D1_O1, Tile_X14Y12_RAM2FAB_D1_O2, Tile_X14Y12_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X14Y12_B (.O0(Tile_X14Y12_RAM2FAB_D1_O0), .O1(Tile_X14Y12_RAM2FAB_D1_O1), .O2(Tile_X14Y12_RAM2FAB_D1_O2), .O3(Tile_X14Y12_RAM2FAB_D1_O3));

wire Tile_X14Y12_RAM2FAB_D2_O0, Tile_X14Y12_RAM2FAB_D2_O1, Tile_X14Y12_RAM2FAB_D2_O2, Tile_X14Y12_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X14Y12_C (.O0(Tile_X14Y12_RAM2FAB_D2_O0), .O1(Tile_X14Y12_RAM2FAB_D2_O1), .O2(Tile_X14Y12_RAM2FAB_D2_O2), .O3(Tile_X14Y12_RAM2FAB_D2_O3));

wire Tile_X14Y12_RAM2FAB_D3_O0, Tile_X14Y12_RAM2FAB_D3_O1, Tile_X14Y12_RAM2FAB_D3_O2, Tile_X14Y12_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X14Y12_D (.O0(Tile_X14Y12_RAM2FAB_D3_O0), .O1(Tile_X14Y12_RAM2FAB_D3_O1), .O2(Tile_X14Y12_RAM2FAB_D3_O2), .O3(Tile_X14Y12_RAM2FAB_D3_O3));

wire Tile_X14Y12_FAB2RAM_D0_I0, Tile_X14Y12_FAB2RAM_D0_I1, Tile_X14Y12_FAB2RAM_D0_I2, Tile_X14Y12_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X14Y12_E (.I0(Tile_X14Y12_FAB2RAM_D0_I0), .I1(Tile_X14Y12_FAB2RAM_D0_I1), .I2(Tile_X14Y12_FAB2RAM_D0_I2), .I3(Tile_X14Y12_FAB2RAM_D0_I3));

wire Tile_X14Y12_FAB2RAM_D1_I0, Tile_X14Y12_FAB2RAM_D1_I1, Tile_X14Y12_FAB2RAM_D1_I2, Tile_X14Y12_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X14Y12_F (.I0(Tile_X14Y12_FAB2RAM_D1_I0), .I1(Tile_X14Y12_FAB2RAM_D1_I1), .I2(Tile_X14Y12_FAB2RAM_D1_I2), .I3(Tile_X14Y12_FAB2RAM_D1_I3));

wire Tile_X14Y12_FAB2RAM_D2_I0, Tile_X14Y12_FAB2RAM_D2_I1, Tile_X14Y12_FAB2RAM_D2_I2, Tile_X14Y12_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X14Y12_G (.I0(Tile_X14Y12_FAB2RAM_D2_I0), .I1(Tile_X14Y12_FAB2RAM_D2_I1), .I2(Tile_X14Y12_FAB2RAM_D2_I2), .I3(Tile_X14Y12_FAB2RAM_D2_I3));

wire Tile_X14Y12_FAB2RAM_D3_I0, Tile_X14Y12_FAB2RAM_D3_I1, Tile_X14Y12_FAB2RAM_D3_I2, Tile_X14Y12_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X14Y12_H (.I0(Tile_X14Y12_FAB2RAM_D3_I0), .I1(Tile_X14Y12_FAB2RAM_D3_I1), .I2(Tile_X14Y12_FAB2RAM_D3_I2), .I3(Tile_X14Y12_FAB2RAM_D3_I3));

wire Tile_X14Y12_FAB2RAM_A0_I0, Tile_X14Y12_FAB2RAM_A0_I1, Tile_X14Y12_FAB2RAM_A0_I2, Tile_X14Y12_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X14Y12_I (.I0(Tile_X14Y12_FAB2RAM_A0_I0), .I1(Tile_X14Y12_FAB2RAM_A0_I1), .I2(Tile_X14Y12_FAB2RAM_A0_I2), .I3(Tile_X14Y12_FAB2RAM_A0_I3));

wire Tile_X14Y12_FAB2RAM_A1_I0, Tile_X14Y12_FAB2RAM_A1_I1, Tile_X14Y12_FAB2RAM_A1_I2, Tile_X14Y12_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X14Y12_J (.I0(Tile_X14Y12_FAB2RAM_A1_I0), .I1(Tile_X14Y12_FAB2RAM_A1_I1), .I2(Tile_X14Y12_FAB2RAM_A1_I2), .I3(Tile_X14Y12_FAB2RAM_A1_I3));

wire Tile_X14Y12_FAB2RAM_C_I0, Tile_X14Y12_FAB2RAM_C_I1, Tile_X14Y12_FAB2RAM_C_I2, Tile_X14Y12_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X14Y12_K (.I0(Tile_X14Y12_FAB2RAM_C_I0), .I1(Tile_X14Y12_FAB2RAM_C_I1), .I2(Tile_X14Y12_FAB2RAM_C_I2), .I3(Tile_X14Y12_FAB2RAM_C_I3));

wire Tile_X0Y13_A_I, Tile_X0Y13_A_T, Tile_X0Y13_A_O, Tile_X0Y13_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y13_A (.O(Tile_X0Y13_A_O), .Q(Tile_X0Y13_A_Q), .I(Tile_X0Y13_A_I));

wire Tile_X0Y13_B_I, Tile_X0Y13_B_T, Tile_X0Y13_B_O, Tile_X0Y13_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y13_B (.O(Tile_X0Y13_B_O), .Q(Tile_X0Y13_B_Q), .I(Tile_X0Y13_B_I));

wire Tile_X14Y13_RAM2FAB_D0_O0, Tile_X14Y13_RAM2FAB_D0_O1, Tile_X14Y13_RAM2FAB_D0_O2, Tile_X14Y13_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X14Y13_A (.O0(Tile_X14Y13_RAM2FAB_D0_O0), .O1(Tile_X14Y13_RAM2FAB_D0_O1), .O2(Tile_X14Y13_RAM2FAB_D0_O2), .O3(Tile_X14Y13_RAM2FAB_D0_O3));

wire Tile_X14Y13_RAM2FAB_D1_O0, Tile_X14Y13_RAM2FAB_D1_O1, Tile_X14Y13_RAM2FAB_D1_O2, Tile_X14Y13_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X14Y13_B (.O0(Tile_X14Y13_RAM2FAB_D1_O0), .O1(Tile_X14Y13_RAM2FAB_D1_O1), .O2(Tile_X14Y13_RAM2FAB_D1_O2), .O3(Tile_X14Y13_RAM2FAB_D1_O3));

wire Tile_X14Y13_RAM2FAB_D2_O0, Tile_X14Y13_RAM2FAB_D2_O1, Tile_X14Y13_RAM2FAB_D2_O2, Tile_X14Y13_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X14Y13_C (.O0(Tile_X14Y13_RAM2FAB_D2_O0), .O1(Tile_X14Y13_RAM2FAB_D2_O1), .O2(Tile_X14Y13_RAM2FAB_D2_O2), .O3(Tile_X14Y13_RAM2FAB_D2_O3));

wire Tile_X14Y13_RAM2FAB_D3_O0, Tile_X14Y13_RAM2FAB_D3_O1, Tile_X14Y13_RAM2FAB_D3_O2, Tile_X14Y13_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X14Y13_D (.O0(Tile_X14Y13_RAM2FAB_D3_O0), .O1(Tile_X14Y13_RAM2FAB_D3_O1), .O2(Tile_X14Y13_RAM2FAB_D3_O2), .O3(Tile_X14Y13_RAM2FAB_D3_O3));

wire Tile_X14Y13_FAB2RAM_D0_I0, Tile_X14Y13_FAB2RAM_D0_I1, Tile_X14Y13_FAB2RAM_D0_I2, Tile_X14Y13_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X14Y13_E (.I0(Tile_X14Y13_FAB2RAM_D0_I0), .I1(Tile_X14Y13_FAB2RAM_D0_I1), .I2(Tile_X14Y13_FAB2RAM_D0_I2), .I3(Tile_X14Y13_FAB2RAM_D0_I3));

wire Tile_X14Y13_FAB2RAM_D1_I0, Tile_X14Y13_FAB2RAM_D1_I1, Tile_X14Y13_FAB2RAM_D1_I2, Tile_X14Y13_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X14Y13_F (.I0(Tile_X14Y13_FAB2RAM_D1_I0), .I1(Tile_X14Y13_FAB2RAM_D1_I1), .I2(Tile_X14Y13_FAB2RAM_D1_I2), .I3(Tile_X14Y13_FAB2RAM_D1_I3));

wire Tile_X14Y13_FAB2RAM_D2_I0, Tile_X14Y13_FAB2RAM_D2_I1, Tile_X14Y13_FAB2RAM_D2_I2, Tile_X14Y13_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X14Y13_G (.I0(Tile_X14Y13_FAB2RAM_D2_I0), .I1(Tile_X14Y13_FAB2RAM_D2_I1), .I2(Tile_X14Y13_FAB2RAM_D2_I2), .I3(Tile_X14Y13_FAB2RAM_D2_I3));

wire Tile_X14Y13_FAB2RAM_D3_I0, Tile_X14Y13_FAB2RAM_D3_I1, Tile_X14Y13_FAB2RAM_D3_I2, Tile_X14Y13_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X14Y13_H (.I0(Tile_X14Y13_FAB2RAM_D3_I0), .I1(Tile_X14Y13_FAB2RAM_D3_I1), .I2(Tile_X14Y13_FAB2RAM_D3_I2), .I3(Tile_X14Y13_FAB2RAM_D3_I3));

wire Tile_X14Y13_FAB2RAM_A0_I0, Tile_X14Y13_FAB2RAM_A0_I1, Tile_X14Y13_FAB2RAM_A0_I2, Tile_X14Y13_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X14Y13_I (.I0(Tile_X14Y13_FAB2RAM_A0_I0), .I1(Tile_X14Y13_FAB2RAM_A0_I1), .I2(Tile_X14Y13_FAB2RAM_A0_I2), .I3(Tile_X14Y13_FAB2RAM_A0_I3));

wire Tile_X14Y13_FAB2RAM_A1_I0, Tile_X14Y13_FAB2RAM_A1_I1, Tile_X14Y13_FAB2RAM_A1_I2, Tile_X14Y13_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X14Y13_J (.I0(Tile_X14Y13_FAB2RAM_A1_I0), .I1(Tile_X14Y13_FAB2RAM_A1_I1), .I2(Tile_X14Y13_FAB2RAM_A1_I2), .I3(Tile_X14Y13_FAB2RAM_A1_I3));

wire Tile_X14Y13_FAB2RAM_C_I0, Tile_X14Y13_FAB2RAM_C_I1, Tile_X14Y13_FAB2RAM_C_I2, Tile_X14Y13_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X14Y13_K (.I0(Tile_X14Y13_FAB2RAM_C_I0), .I1(Tile_X14Y13_FAB2RAM_C_I1), .I2(Tile_X14Y13_FAB2RAM_C_I2), .I3(Tile_X14Y13_FAB2RAM_C_I3));

wire Tile_X0Y14_A_I, Tile_X0Y14_A_T, Tile_X0Y14_A_O, Tile_X0Y14_A_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y14_A (.O(Tile_X0Y14_A_O), .Q(Tile_X0Y14_A_Q), .I(Tile_X0Y14_A_I));

wire Tile_X0Y14_B_I, Tile_X0Y14_B_T, Tile_X0Y14_B_O, Tile_X0Y14_B_Q;
(* keep *) IO_1_bidirectional_frame_config_pass Tile_X0Y14_B (.O(Tile_X0Y14_B_O), .Q(Tile_X0Y14_B_Q), .I(Tile_X0Y14_B_I));

wire Tile_X14Y14_RAM2FAB_D0_O0, Tile_X14Y14_RAM2FAB_D0_O1, Tile_X14Y14_RAM2FAB_D0_O2, Tile_X14Y14_RAM2FAB_D0_O3;
(* keep *) InPass4_frame_config Tile_X14Y14_A (.O0(Tile_X14Y14_RAM2FAB_D0_O0), .O1(Tile_X14Y14_RAM2FAB_D0_O1), .O2(Tile_X14Y14_RAM2FAB_D0_O2), .O3(Tile_X14Y14_RAM2FAB_D0_O3));

wire Tile_X14Y14_RAM2FAB_D1_O0, Tile_X14Y14_RAM2FAB_D1_O1, Tile_X14Y14_RAM2FAB_D1_O2, Tile_X14Y14_RAM2FAB_D1_O3;
(* keep *) InPass4_frame_config Tile_X14Y14_B (.O0(Tile_X14Y14_RAM2FAB_D1_O0), .O1(Tile_X14Y14_RAM2FAB_D1_O1), .O2(Tile_X14Y14_RAM2FAB_D1_O2), .O3(Tile_X14Y14_RAM2FAB_D1_O3));

wire Tile_X14Y14_RAM2FAB_D2_O0, Tile_X14Y14_RAM2FAB_D2_O1, Tile_X14Y14_RAM2FAB_D2_O2, Tile_X14Y14_RAM2FAB_D2_O3;
(* keep *) InPass4_frame_config Tile_X14Y14_C (.O0(Tile_X14Y14_RAM2FAB_D2_O0), .O1(Tile_X14Y14_RAM2FAB_D2_O1), .O2(Tile_X14Y14_RAM2FAB_D2_O2), .O3(Tile_X14Y14_RAM2FAB_D2_O3));

wire Tile_X14Y14_RAM2FAB_D3_O0, Tile_X14Y14_RAM2FAB_D3_O1, Tile_X14Y14_RAM2FAB_D3_O2, Tile_X14Y14_RAM2FAB_D3_O3;
(* keep *) InPass4_frame_config Tile_X14Y14_D (.O0(Tile_X14Y14_RAM2FAB_D3_O0), .O1(Tile_X14Y14_RAM2FAB_D3_O1), .O2(Tile_X14Y14_RAM2FAB_D3_O2), .O3(Tile_X14Y14_RAM2FAB_D3_O3));

wire Tile_X14Y14_FAB2RAM_D0_I0, Tile_X14Y14_FAB2RAM_D0_I1, Tile_X14Y14_FAB2RAM_D0_I2, Tile_X14Y14_FAB2RAM_D0_I3;
(* keep *) OutPass4_frame_config Tile_X14Y14_E (.I0(Tile_X14Y14_FAB2RAM_D0_I0), .I1(Tile_X14Y14_FAB2RAM_D0_I1), .I2(Tile_X14Y14_FAB2RAM_D0_I2), .I3(Tile_X14Y14_FAB2RAM_D0_I3));

wire Tile_X14Y14_FAB2RAM_D1_I0, Tile_X14Y14_FAB2RAM_D1_I1, Tile_X14Y14_FAB2RAM_D1_I2, Tile_X14Y14_FAB2RAM_D1_I3;
(* keep *) OutPass4_frame_config Tile_X14Y14_F (.I0(Tile_X14Y14_FAB2RAM_D1_I0), .I1(Tile_X14Y14_FAB2RAM_D1_I1), .I2(Tile_X14Y14_FAB2RAM_D1_I2), .I3(Tile_X14Y14_FAB2RAM_D1_I3));

wire Tile_X14Y14_FAB2RAM_D2_I0, Tile_X14Y14_FAB2RAM_D2_I1, Tile_X14Y14_FAB2RAM_D2_I2, Tile_X14Y14_FAB2RAM_D2_I3;
(* keep *) OutPass4_frame_config Tile_X14Y14_G (.I0(Tile_X14Y14_FAB2RAM_D2_I0), .I1(Tile_X14Y14_FAB2RAM_D2_I1), .I2(Tile_X14Y14_FAB2RAM_D2_I2), .I3(Tile_X14Y14_FAB2RAM_D2_I3));

wire Tile_X14Y14_FAB2RAM_D3_I0, Tile_X14Y14_FAB2RAM_D3_I1, Tile_X14Y14_FAB2RAM_D3_I2, Tile_X14Y14_FAB2RAM_D3_I3;
(* keep *) OutPass4_frame_config Tile_X14Y14_H (.I0(Tile_X14Y14_FAB2RAM_D3_I0), .I1(Tile_X14Y14_FAB2RAM_D3_I1), .I2(Tile_X14Y14_FAB2RAM_D3_I2), .I3(Tile_X14Y14_FAB2RAM_D3_I3));

wire Tile_X14Y14_FAB2RAM_A0_I0, Tile_X14Y14_FAB2RAM_A0_I1, Tile_X14Y14_FAB2RAM_A0_I2, Tile_X14Y14_FAB2RAM_A0_I3;
(* keep *) OutPass4_frame_config Tile_X14Y14_I (.I0(Tile_X14Y14_FAB2RAM_A0_I0), .I1(Tile_X14Y14_FAB2RAM_A0_I1), .I2(Tile_X14Y14_FAB2RAM_A0_I2), .I3(Tile_X14Y14_FAB2RAM_A0_I3));

wire Tile_X14Y14_FAB2RAM_A1_I0, Tile_X14Y14_FAB2RAM_A1_I1, Tile_X14Y14_FAB2RAM_A1_I2, Tile_X14Y14_FAB2RAM_A1_I3;
(* keep *) OutPass4_frame_config Tile_X14Y14_J (.I0(Tile_X14Y14_FAB2RAM_A1_I0), .I1(Tile_X14Y14_FAB2RAM_A1_I1), .I2(Tile_X14Y14_FAB2RAM_A1_I2), .I3(Tile_X14Y14_FAB2RAM_A1_I3));

wire Tile_X14Y14_FAB2RAM_C_I0, Tile_X14Y14_FAB2RAM_C_I1, Tile_X14Y14_FAB2RAM_C_I2, Tile_X14Y14_FAB2RAM_C_I3;
(* keep *) OutPass4_frame_config Tile_X14Y14_K (.I0(Tile_X14Y14_FAB2RAM_C_I0), .I1(Tile_X14Y14_FAB2RAM_C_I1), .I2(Tile_X14Y14_FAB2RAM_C_I2), .I3(Tile_X14Y14_FAB2RAM_C_I3));

endmodule